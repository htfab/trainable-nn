magic
tech sky130B
magscale 1 2
timestamp 1663010149
<< obsli1 >>
rect 1104 2159 358892 477649
<< obsm1 >>
rect 290 280 358892 477680
<< metal2 >>
rect 3238 479200 3294 480000
rect 6366 479200 6422 480000
rect 9494 479200 9550 480000
rect 12622 479200 12678 480000
rect 15750 479200 15806 480000
rect 18878 479200 18934 480000
rect 22006 479200 22062 480000
rect 25134 479200 25190 480000
rect 28262 479200 28318 480000
rect 31390 479200 31446 480000
rect 34518 479200 34574 480000
rect 37646 479200 37702 480000
rect 40774 479200 40830 480000
rect 43902 479200 43958 480000
rect 47030 479200 47086 480000
rect 50158 479200 50214 480000
rect 53286 479200 53342 480000
rect 56414 479200 56470 480000
rect 59542 479200 59598 480000
rect 62670 479200 62726 480000
rect 65798 479200 65854 480000
rect 68926 479200 68982 480000
rect 72054 479200 72110 480000
rect 75182 479200 75238 480000
rect 78310 479200 78366 480000
rect 81438 479200 81494 480000
rect 84566 479200 84622 480000
rect 87694 479200 87750 480000
rect 90822 479200 90878 480000
rect 93950 479200 94006 480000
rect 97078 479200 97134 480000
rect 100206 479200 100262 480000
rect 103334 479200 103390 480000
rect 106462 479200 106518 480000
rect 109590 479200 109646 480000
rect 112718 479200 112774 480000
rect 115846 479200 115902 480000
rect 118974 479200 119030 480000
rect 122102 479200 122158 480000
rect 125230 479200 125286 480000
rect 128358 479200 128414 480000
rect 131486 479200 131542 480000
rect 134614 479200 134670 480000
rect 137742 479200 137798 480000
rect 140870 479200 140926 480000
rect 143998 479200 144054 480000
rect 147126 479200 147182 480000
rect 150254 479200 150310 480000
rect 153382 479200 153438 480000
rect 156510 479200 156566 480000
rect 159638 479200 159694 480000
rect 162766 479200 162822 480000
rect 165894 479200 165950 480000
rect 169022 479200 169078 480000
rect 172150 479200 172206 480000
rect 175278 479200 175334 480000
rect 178406 479200 178462 480000
rect 181534 479200 181590 480000
rect 184662 479200 184718 480000
rect 187790 479200 187846 480000
rect 190918 479200 190974 480000
rect 194046 479200 194102 480000
rect 197174 479200 197230 480000
rect 200302 479200 200358 480000
rect 203430 479200 203486 480000
rect 206558 479200 206614 480000
rect 209686 479200 209742 480000
rect 212814 479200 212870 480000
rect 215942 479200 215998 480000
rect 219070 479200 219126 480000
rect 222198 479200 222254 480000
rect 225326 479200 225382 480000
rect 228454 479200 228510 480000
rect 231582 479200 231638 480000
rect 234710 479200 234766 480000
rect 237838 479200 237894 480000
rect 240966 479200 241022 480000
rect 244094 479200 244150 480000
rect 247222 479200 247278 480000
rect 250350 479200 250406 480000
rect 253478 479200 253534 480000
rect 256606 479200 256662 480000
rect 259734 479200 259790 480000
rect 262862 479200 262918 480000
rect 265990 479200 266046 480000
rect 269118 479200 269174 480000
rect 272246 479200 272302 480000
rect 275374 479200 275430 480000
rect 278502 479200 278558 480000
rect 281630 479200 281686 480000
rect 284758 479200 284814 480000
rect 287886 479200 287942 480000
rect 291014 479200 291070 480000
rect 294142 479200 294198 480000
rect 297270 479200 297326 480000
rect 300398 479200 300454 480000
rect 303526 479200 303582 480000
rect 306654 479200 306710 480000
rect 309782 479200 309838 480000
rect 312910 479200 312966 480000
rect 316038 479200 316094 480000
rect 319166 479200 319222 480000
rect 322294 479200 322350 480000
rect 325422 479200 325478 480000
rect 328550 479200 328606 480000
rect 331678 479200 331734 480000
rect 334806 479200 334862 480000
rect 337934 479200 337990 480000
rect 341062 479200 341118 480000
rect 344190 479200 344246 480000
rect 347318 479200 347374 480000
rect 350446 479200 350502 480000
rect 353574 479200 353630 480000
rect 356702 479200 356758 480000
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22834 0 22890 800
rect 23478 0 23534 800
rect 24122 0 24178 800
rect 24766 0 24822 800
rect 25410 0 25466 800
rect 26054 0 26110 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29274 0 29330 800
rect 29918 0 29974 800
rect 30562 0 30618 800
rect 31206 0 31262 800
rect 31850 0 31906 800
rect 32494 0 32550 800
rect 33138 0 33194 800
rect 33782 0 33838 800
rect 34426 0 34482 800
rect 35070 0 35126 800
rect 35714 0 35770 800
rect 36358 0 36414 800
rect 37002 0 37058 800
rect 37646 0 37702 800
rect 38290 0 38346 800
rect 38934 0 38990 800
rect 39578 0 39634 800
rect 40222 0 40278 800
rect 40866 0 40922 800
rect 41510 0 41566 800
rect 42154 0 42210 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 44086 0 44142 800
rect 44730 0 44786 800
rect 45374 0 45430 800
rect 46018 0 46074 800
rect 46662 0 46718 800
rect 47306 0 47362 800
rect 47950 0 48006 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55678 0 55734 800
rect 56322 0 56378 800
rect 56966 0 57022 800
rect 57610 0 57666 800
rect 58254 0 58310 800
rect 58898 0 58954 800
rect 59542 0 59598 800
rect 60186 0 60242 800
rect 60830 0 60886 800
rect 61474 0 61530 800
rect 62118 0 62174 800
rect 62762 0 62818 800
rect 63406 0 63462 800
rect 64050 0 64106 800
rect 64694 0 64750 800
rect 65338 0 65394 800
rect 65982 0 66038 800
rect 66626 0 66682 800
rect 67270 0 67326 800
rect 67914 0 67970 800
rect 68558 0 68614 800
rect 69202 0 69258 800
rect 69846 0 69902 800
rect 70490 0 70546 800
rect 71134 0 71190 800
rect 71778 0 71834 800
rect 72422 0 72478 800
rect 73066 0 73122 800
rect 73710 0 73766 800
rect 74354 0 74410 800
rect 74998 0 75054 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 76930 0 76986 800
rect 77574 0 77630 800
rect 78218 0 78274 800
rect 78862 0 78918 800
rect 79506 0 79562 800
rect 80150 0 80206 800
rect 80794 0 80850 800
rect 81438 0 81494 800
rect 82082 0 82138 800
rect 82726 0 82782 800
rect 83370 0 83426 800
rect 84014 0 84070 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 85946 0 86002 800
rect 86590 0 86646 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89166 0 89222 800
rect 89810 0 89866 800
rect 90454 0 90510 800
rect 91098 0 91154 800
rect 91742 0 91798 800
rect 92386 0 92442 800
rect 93030 0 93086 800
rect 93674 0 93730 800
rect 94318 0 94374 800
rect 94962 0 95018 800
rect 95606 0 95662 800
rect 96250 0 96306 800
rect 96894 0 96950 800
rect 97538 0 97594 800
rect 98182 0 98238 800
rect 98826 0 98882 800
rect 99470 0 99526 800
rect 100114 0 100170 800
rect 100758 0 100814 800
rect 101402 0 101458 800
rect 102046 0 102102 800
rect 102690 0 102746 800
rect 103334 0 103390 800
rect 103978 0 104034 800
rect 104622 0 104678 800
rect 105266 0 105322 800
rect 105910 0 105966 800
rect 106554 0 106610 800
rect 107198 0 107254 800
rect 107842 0 107898 800
rect 108486 0 108542 800
rect 109130 0 109186 800
rect 109774 0 109830 800
rect 110418 0 110474 800
rect 111062 0 111118 800
rect 111706 0 111762 800
rect 112350 0 112406 800
rect 112994 0 113050 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114926 0 114982 800
rect 115570 0 115626 800
rect 116214 0 116270 800
rect 116858 0 116914 800
rect 117502 0 117558 800
rect 118146 0 118202 800
rect 118790 0 118846 800
rect 119434 0 119490 800
rect 120078 0 120134 800
rect 120722 0 120778 800
rect 121366 0 121422 800
rect 122010 0 122066 800
rect 122654 0 122710 800
rect 123298 0 123354 800
rect 123942 0 123998 800
rect 124586 0 124642 800
rect 125230 0 125286 800
rect 125874 0 125930 800
rect 126518 0 126574 800
rect 127162 0 127218 800
rect 127806 0 127862 800
rect 128450 0 128506 800
rect 129094 0 129150 800
rect 129738 0 129794 800
rect 130382 0 130438 800
rect 131026 0 131082 800
rect 131670 0 131726 800
rect 132314 0 132370 800
rect 132958 0 133014 800
rect 133602 0 133658 800
rect 134246 0 134302 800
rect 134890 0 134946 800
rect 135534 0 135590 800
rect 136178 0 136234 800
rect 136822 0 136878 800
rect 137466 0 137522 800
rect 138110 0 138166 800
rect 138754 0 138810 800
rect 139398 0 139454 800
rect 140042 0 140098 800
rect 140686 0 140742 800
rect 141330 0 141386 800
rect 141974 0 142030 800
rect 142618 0 142674 800
rect 143262 0 143318 800
rect 143906 0 143962 800
rect 144550 0 144606 800
rect 145194 0 145250 800
rect 145838 0 145894 800
rect 146482 0 146538 800
rect 147126 0 147182 800
rect 147770 0 147826 800
rect 148414 0 148470 800
rect 149058 0 149114 800
rect 149702 0 149758 800
rect 150346 0 150402 800
rect 150990 0 151046 800
rect 151634 0 151690 800
rect 152278 0 152334 800
rect 152922 0 152978 800
rect 153566 0 153622 800
rect 154210 0 154266 800
rect 154854 0 154910 800
rect 155498 0 155554 800
rect 156142 0 156198 800
rect 156786 0 156842 800
rect 157430 0 157486 800
rect 158074 0 158130 800
rect 158718 0 158774 800
rect 159362 0 159418 800
rect 160006 0 160062 800
rect 160650 0 160706 800
rect 161294 0 161350 800
rect 161938 0 161994 800
rect 162582 0 162638 800
rect 163226 0 163282 800
rect 163870 0 163926 800
rect 164514 0 164570 800
rect 165158 0 165214 800
rect 165802 0 165858 800
rect 166446 0 166502 800
rect 167090 0 167146 800
rect 167734 0 167790 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169666 0 169722 800
rect 170310 0 170366 800
rect 170954 0 171010 800
rect 171598 0 171654 800
rect 172242 0 172298 800
rect 172886 0 172942 800
rect 173530 0 173586 800
rect 174174 0 174230 800
rect 174818 0 174874 800
rect 175462 0 175518 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177394 0 177450 800
rect 178038 0 178094 800
rect 178682 0 178738 800
rect 179326 0 179382 800
rect 179970 0 180026 800
rect 180614 0 180670 800
rect 181258 0 181314 800
rect 181902 0 181958 800
rect 182546 0 182602 800
rect 183190 0 183246 800
rect 183834 0 183890 800
rect 184478 0 184534 800
rect 185122 0 185178 800
rect 185766 0 185822 800
rect 186410 0 186466 800
rect 187054 0 187110 800
rect 187698 0 187754 800
rect 188342 0 188398 800
rect 188986 0 189042 800
rect 189630 0 189686 800
rect 190274 0 190330 800
rect 190918 0 190974 800
rect 191562 0 191618 800
rect 192206 0 192262 800
rect 192850 0 192906 800
rect 193494 0 193550 800
rect 194138 0 194194 800
rect 194782 0 194838 800
rect 195426 0 195482 800
rect 196070 0 196126 800
rect 196714 0 196770 800
rect 197358 0 197414 800
rect 198002 0 198058 800
rect 198646 0 198702 800
rect 199290 0 199346 800
rect 199934 0 199990 800
rect 200578 0 200634 800
rect 201222 0 201278 800
rect 201866 0 201922 800
rect 202510 0 202566 800
rect 203154 0 203210 800
rect 203798 0 203854 800
rect 204442 0 204498 800
rect 205086 0 205142 800
rect 205730 0 205786 800
rect 206374 0 206430 800
rect 207018 0 207074 800
rect 207662 0 207718 800
rect 208306 0 208362 800
rect 208950 0 209006 800
rect 209594 0 209650 800
rect 210238 0 210294 800
rect 210882 0 210938 800
rect 211526 0 211582 800
rect 212170 0 212226 800
rect 212814 0 212870 800
rect 213458 0 213514 800
rect 214102 0 214158 800
rect 214746 0 214802 800
rect 215390 0 215446 800
rect 216034 0 216090 800
rect 216678 0 216734 800
rect 217322 0 217378 800
rect 217966 0 218022 800
rect 218610 0 218666 800
rect 219254 0 219310 800
rect 219898 0 219954 800
rect 220542 0 220598 800
rect 221186 0 221242 800
rect 221830 0 221886 800
rect 222474 0 222530 800
rect 223118 0 223174 800
rect 223762 0 223818 800
rect 224406 0 224462 800
rect 225050 0 225106 800
rect 225694 0 225750 800
rect 226338 0 226394 800
rect 226982 0 227038 800
rect 227626 0 227682 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229558 0 229614 800
rect 230202 0 230258 800
rect 230846 0 230902 800
rect 231490 0 231546 800
rect 232134 0 232190 800
rect 232778 0 232834 800
rect 233422 0 233478 800
rect 234066 0 234122 800
rect 234710 0 234766 800
rect 235354 0 235410 800
rect 235998 0 236054 800
rect 236642 0 236698 800
rect 237286 0 237342 800
rect 237930 0 237986 800
rect 238574 0 238630 800
rect 239218 0 239274 800
rect 239862 0 239918 800
rect 240506 0 240562 800
rect 241150 0 241206 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 243082 0 243138 800
rect 243726 0 243782 800
rect 244370 0 244426 800
rect 245014 0 245070 800
rect 245658 0 245714 800
rect 246302 0 246358 800
rect 246946 0 247002 800
rect 247590 0 247646 800
rect 248234 0 248290 800
rect 248878 0 248934 800
rect 249522 0 249578 800
rect 250166 0 250222 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252098 0 252154 800
rect 252742 0 252798 800
rect 253386 0 253442 800
rect 254030 0 254086 800
rect 254674 0 254730 800
rect 255318 0 255374 800
rect 255962 0 256018 800
rect 256606 0 256662 800
rect 257250 0 257306 800
rect 257894 0 257950 800
rect 258538 0 258594 800
rect 259182 0 259238 800
rect 259826 0 259882 800
rect 260470 0 260526 800
rect 261114 0 261170 800
rect 261758 0 261814 800
rect 262402 0 262458 800
rect 263046 0 263102 800
rect 263690 0 263746 800
rect 264334 0 264390 800
rect 264978 0 265034 800
rect 265622 0 265678 800
rect 266266 0 266322 800
rect 266910 0 266966 800
rect 267554 0 267610 800
rect 268198 0 268254 800
rect 268842 0 268898 800
rect 269486 0 269542 800
rect 270130 0 270186 800
rect 270774 0 270830 800
rect 271418 0 271474 800
rect 272062 0 272118 800
rect 272706 0 272762 800
rect 273350 0 273406 800
rect 273994 0 274050 800
rect 274638 0 274694 800
rect 275282 0 275338 800
rect 275926 0 275982 800
rect 276570 0 276626 800
rect 277214 0 277270 800
rect 277858 0 277914 800
rect 278502 0 278558 800
rect 279146 0 279202 800
rect 279790 0 279846 800
rect 280434 0 280490 800
rect 281078 0 281134 800
rect 281722 0 281778 800
rect 282366 0 282422 800
rect 283010 0 283066 800
rect 283654 0 283710 800
rect 284298 0 284354 800
rect 284942 0 284998 800
rect 285586 0 285642 800
rect 286230 0 286286 800
rect 286874 0 286930 800
rect 287518 0 287574 800
rect 288162 0 288218 800
rect 288806 0 288862 800
rect 289450 0 289506 800
rect 290094 0 290150 800
rect 290738 0 290794 800
rect 291382 0 291438 800
rect 292026 0 292082 800
rect 292670 0 292726 800
rect 293314 0 293370 800
rect 293958 0 294014 800
rect 294602 0 294658 800
rect 295246 0 295302 800
rect 295890 0 295946 800
rect 296534 0 296590 800
rect 297178 0 297234 800
rect 297822 0 297878 800
rect 298466 0 298522 800
rect 299110 0 299166 800
rect 299754 0 299810 800
rect 300398 0 300454 800
rect 301042 0 301098 800
rect 301686 0 301742 800
rect 302330 0 302386 800
rect 302974 0 303030 800
rect 303618 0 303674 800
rect 304262 0 304318 800
rect 304906 0 304962 800
rect 305550 0 305606 800
rect 306194 0 306250 800
rect 306838 0 306894 800
rect 307482 0 307538 800
rect 308126 0 308182 800
rect 308770 0 308826 800
rect 309414 0 309470 800
rect 310058 0 310114 800
rect 310702 0 310758 800
rect 311346 0 311402 800
rect 311990 0 312046 800
rect 312634 0 312690 800
rect 313278 0 313334 800
rect 313922 0 313978 800
rect 314566 0 314622 800
rect 315210 0 315266 800
rect 315854 0 315910 800
rect 316498 0 316554 800
rect 317142 0 317198 800
rect 317786 0 317842 800
rect 318430 0 318486 800
rect 319074 0 319130 800
rect 319718 0 319774 800
rect 320362 0 320418 800
rect 321006 0 321062 800
rect 321650 0 321706 800
rect 322294 0 322350 800
rect 322938 0 322994 800
rect 323582 0 323638 800
rect 324226 0 324282 800
rect 324870 0 324926 800
rect 325514 0 325570 800
rect 326158 0 326214 800
rect 326802 0 326858 800
rect 327446 0 327502 800
rect 328090 0 328146 800
rect 328734 0 328790 800
rect 329378 0 329434 800
rect 330022 0 330078 800
rect 330666 0 330722 800
rect 331310 0 331366 800
rect 331954 0 332010 800
rect 332598 0 332654 800
rect 333242 0 333298 800
rect 333886 0 333942 800
rect 334530 0 334586 800
rect 335174 0 335230 800
rect 335818 0 335874 800
rect 336462 0 336518 800
rect 337106 0 337162 800
rect 337750 0 337806 800
rect 338394 0 338450 800
<< obsm2 >>
rect 296 479144 3182 479346
rect 3350 479144 6310 479346
rect 6478 479144 9438 479346
rect 9606 479144 12566 479346
rect 12734 479144 15694 479346
rect 15862 479144 18822 479346
rect 18990 479144 21950 479346
rect 22118 479144 25078 479346
rect 25246 479144 28206 479346
rect 28374 479144 31334 479346
rect 31502 479144 34462 479346
rect 34630 479144 37590 479346
rect 37758 479144 40718 479346
rect 40886 479144 43846 479346
rect 44014 479144 46974 479346
rect 47142 479144 50102 479346
rect 50270 479144 53230 479346
rect 53398 479144 56358 479346
rect 56526 479144 59486 479346
rect 59654 479144 62614 479346
rect 62782 479144 65742 479346
rect 65910 479144 68870 479346
rect 69038 479144 71998 479346
rect 72166 479144 75126 479346
rect 75294 479144 78254 479346
rect 78422 479144 81382 479346
rect 81550 479144 84510 479346
rect 84678 479144 87638 479346
rect 87806 479144 90766 479346
rect 90934 479144 93894 479346
rect 94062 479144 97022 479346
rect 97190 479144 100150 479346
rect 100318 479144 103278 479346
rect 103446 479144 106406 479346
rect 106574 479144 109534 479346
rect 109702 479144 112662 479346
rect 112830 479144 115790 479346
rect 115958 479144 118918 479346
rect 119086 479144 122046 479346
rect 122214 479144 125174 479346
rect 125342 479144 128302 479346
rect 128470 479144 131430 479346
rect 131598 479144 134558 479346
rect 134726 479144 137686 479346
rect 137854 479144 140814 479346
rect 140982 479144 143942 479346
rect 144110 479144 147070 479346
rect 147238 479144 150198 479346
rect 150366 479144 153326 479346
rect 153494 479144 156454 479346
rect 156622 479144 159582 479346
rect 159750 479144 162710 479346
rect 162878 479144 165838 479346
rect 166006 479144 168966 479346
rect 169134 479144 172094 479346
rect 172262 479144 175222 479346
rect 175390 479144 178350 479346
rect 178518 479144 181478 479346
rect 181646 479144 184606 479346
rect 184774 479144 187734 479346
rect 187902 479144 190862 479346
rect 191030 479144 193990 479346
rect 194158 479144 197118 479346
rect 197286 479144 200246 479346
rect 200414 479144 203374 479346
rect 203542 479144 206502 479346
rect 206670 479144 209630 479346
rect 209798 479144 212758 479346
rect 212926 479144 215886 479346
rect 216054 479144 219014 479346
rect 219182 479144 222142 479346
rect 222310 479144 225270 479346
rect 225438 479144 228398 479346
rect 228566 479144 231526 479346
rect 231694 479144 234654 479346
rect 234822 479144 237782 479346
rect 237950 479144 240910 479346
rect 241078 479144 244038 479346
rect 244206 479144 247166 479346
rect 247334 479144 250294 479346
rect 250462 479144 253422 479346
rect 253590 479144 256550 479346
rect 256718 479144 259678 479346
rect 259846 479144 262806 479346
rect 262974 479144 265934 479346
rect 266102 479144 269062 479346
rect 269230 479144 272190 479346
rect 272358 479144 275318 479346
rect 275486 479144 278446 479346
rect 278614 479144 281574 479346
rect 281742 479144 284702 479346
rect 284870 479144 287830 479346
rect 287998 479144 290958 479346
rect 291126 479144 294086 479346
rect 294254 479144 297214 479346
rect 297382 479144 300342 479346
rect 300510 479144 303470 479346
rect 303638 479144 306598 479346
rect 306766 479144 309726 479346
rect 309894 479144 312854 479346
rect 313022 479144 315982 479346
rect 316150 479144 319110 479346
rect 319278 479144 322238 479346
rect 322406 479144 325366 479346
rect 325534 479144 328494 479346
rect 328662 479144 331622 479346
rect 331790 479144 334750 479346
rect 334918 479144 337878 479346
rect 338046 479144 341006 479346
rect 341174 479144 344134 479346
rect 344302 479144 347262 479346
rect 347430 479144 350390 479346
rect 350558 479144 353518 479346
rect 353686 479144 356646 479346
rect 356814 479144 358596 479346
rect 296 856 358596 479144
rect 296 274 21490 856
rect 21658 274 22134 856
rect 22302 274 22778 856
rect 22946 274 23422 856
rect 23590 274 24066 856
rect 24234 274 24710 856
rect 24878 274 25354 856
rect 25522 274 25998 856
rect 26166 274 26642 856
rect 26810 274 27286 856
rect 27454 274 27930 856
rect 28098 274 28574 856
rect 28742 274 29218 856
rect 29386 274 29862 856
rect 30030 274 30506 856
rect 30674 274 31150 856
rect 31318 274 31794 856
rect 31962 274 32438 856
rect 32606 274 33082 856
rect 33250 274 33726 856
rect 33894 274 34370 856
rect 34538 274 35014 856
rect 35182 274 35658 856
rect 35826 274 36302 856
rect 36470 274 36946 856
rect 37114 274 37590 856
rect 37758 274 38234 856
rect 38402 274 38878 856
rect 39046 274 39522 856
rect 39690 274 40166 856
rect 40334 274 40810 856
rect 40978 274 41454 856
rect 41622 274 42098 856
rect 42266 274 42742 856
rect 42910 274 43386 856
rect 43554 274 44030 856
rect 44198 274 44674 856
rect 44842 274 45318 856
rect 45486 274 45962 856
rect 46130 274 46606 856
rect 46774 274 47250 856
rect 47418 274 47894 856
rect 48062 274 48538 856
rect 48706 274 49182 856
rect 49350 274 49826 856
rect 49994 274 50470 856
rect 50638 274 51114 856
rect 51282 274 51758 856
rect 51926 274 52402 856
rect 52570 274 53046 856
rect 53214 274 53690 856
rect 53858 274 54334 856
rect 54502 274 54978 856
rect 55146 274 55622 856
rect 55790 274 56266 856
rect 56434 274 56910 856
rect 57078 274 57554 856
rect 57722 274 58198 856
rect 58366 274 58842 856
rect 59010 274 59486 856
rect 59654 274 60130 856
rect 60298 274 60774 856
rect 60942 274 61418 856
rect 61586 274 62062 856
rect 62230 274 62706 856
rect 62874 274 63350 856
rect 63518 274 63994 856
rect 64162 274 64638 856
rect 64806 274 65282 856
rect 65450 274 65926 856
rect 66094 274 66570 856
rect 66738 274 67214 856
rect 67382 274 67858 856
rect 68026 274 68502 856
rect 68670 274 69146 856
rect 69314 274 69790 856
rect 69958 274 70434 856
rect 70602 274 71078 856
rect 71246 274 71722 856
rect 71890 274 72366 856
rect 72534 274 73010 856
rect 73178 274 73654 856
rect 73822 274 74298 856
rect 74466 274 74942 856
rect 75110 274 75586 856
rect 75754 274 76230 856
rect 76398 274 76874 856
rect 77042 274 77518 856
rect 77686 274 78162 856
rect 78330 274 78806 856
rect 78974 274 79450 856
rect 79618 274 80094 856
rect 80262 274 80738 856
rect 80906 274 81382 856
rect 81550 274 82026 856
rect 82194 274 82670 856
rect 82838 274 83314 856
rect 83482 274 83958 856
rect 84126 274 84602 856
rect 84770 274 85246 856
rect 85414 274 85890 856
rect 86058 274 86534 856
rect 86702 274 87178 856
rect 87346 274 87822 856
rect 87990 274 88466 856
rect 88634 274 89110 856
rect 89278 274 89754 856
rect 89922 274 90398 856
rect 90566 274 91042 856
rect 91210 274 91686 856
rect 91854 274 92330 856
rect 92498 274 92974 856
rect 93142 274 93618 856
rect 93786 274 94262 856
rect 94430 274 94906 856
rect 95074 274 95550 856
rect 95718 274 96194 856
rect 96362 274 96838 856
rect 97006 274 97482 856
rect 97650 274 98126 856
rect 98294 274 98770 856
rect 98938 274 99414 856
rect 99582 274 100058 856
rect 100226 274 100702 856
rect 100870 274 101346 856
rect 101514 274 101990 856
rect 102158 274 102634 856
rect 102802 274 103278 856
rect 103446 274 103922 856
rect 104090 274 104566 856
rect 104734 274 105210 856
rect 105378 274 105854 856
rect 106022 274 106498 856
rect 106666 274 107142 856
rect 107310 274 107786 856
rect 107954 274 108430 856
rect 108598 274 109074 856
rect 109242 274 109718 856
rect 109886 274 110362 856
rect 110530 274 111006 856
rect 111174 274 111650 856
rect 111818 274 112294 856
rect 112462 274 112938 856
rect 113106 274 113582 856
rect 113750 274 114226 856
rect 114394 274 114870 856
rect 115038 274 115514 856
rect 115682 274 116158 856
rect 116326 274 116802 856
rect 116970 274 117446 856
rect 117614 274 118090 856
rect 118258 274 118734 856
rect 118902 274 119378 856
rect 119546 274 120022 856
rect 120190 274 120666 856
rect 120834 274 121310 856
rect 121478 274 121954 856
rect 122122 274 122598 856
rect 122766 274 123242 856
rect 123410 274 123886 856
rect 124054 274 124530 856
rect 124698 274 125174 856
rect 125342 274 125818 856
rect 125986 274 126462 856
rect 126630 274 127106 856
rect 127274 274 127750 856
rect 127918 274 128394 856
rect 128562 274 129038 856
rect 129206 274 129682 856
rect 129850 274 130326 856
rect 130494 274 130970 856
rect 131138 274 131614 856
rect 131782 274 132258 856
rect 132426 274 132902 856
rect 133070 274 133546 856
rect 133714 274 134190 856
rect 134358 274 134834 856
rect 135002 274 135478 856
rect 135646 274 136122 856
rect 136290 274 136766 856
rect 136934 274 137410 856
rect 137578 274 138054 856
rect 138222 274 138698 856
rect 138866 274 139342 856
rect 139510 274 139986 856
rect 140154 274 140630 856
rect 140798 274 141274 856
rect 141442 274 141918 856
rect 142086 274 142562 856
rect 142730 274 143206 856
rect 143374 274 143850 856
rect 144018 274 144494 856
rect 144662 274 145138 856
rect 145306 274 145782 856
rect 145950 274 146426 856
rect 146594 274 147070 856
rect 147238 274 147714 856
rect 147882 274 148358 856
rect 148526 274 149002 856
rect 149170 274 149646 856
rect 149814 274 150290 856
rect 150458 274 150934 856
rect 151102 274 151578 856
rect 151746 274 152222 856
rect 152390 274 152866 856
rect 153034 274 153510 856
rect 153678 274 154154 856
rect 154322 274 154798 856
rect 154966 274 155442 856
rect 155610 274 156086 856
rect 156254 274 156730 856
rect 156898 274 157374 856
rect 157542 274 158018 856
rect 158186 274 158662 856
rect 158830 274 159306 856
rect 159474 274 159950 856
rect 160118 274 160594 856
rect 160762 274 161238 856
rect 161406 274 161882 856
rect 162050 274 162526 856
rect 162694 274 163170 856
rect 163338 274 163814 856
rect 163982 274 164458 856
rect 164626 274 165102 856
rect 165270 274 165746 856
rect 165914 274 166390 856
rect 166558 274 167034 856
rect 167202 274 167678 856
rect 167846 274 168322 856
rect 168490 274 168966 856
rect 169134 274 169610 856
rect 169778 274 170254 856
rect 170422 274 170898 856
rect 171066 274 171542 856
rect 171710 274 172186 856
rect 172354 274 172830 856
rect 172998 274 173474 856
rect 173642 274 174118 856
rect 174286 274 174762 856
rect 174930 274 175406 856
rect 175574 274 176050 856
rect 176218 274 176694 856
rect 176862 274 177338 856
rect 177506 274 177982 856
rect 178150 274 178626 856
rect 178794 274 179270 856
rect 179438 274 179914 856
rect 180082 274 180558 856
rect 180726 274 181202 856
rect 181370 274 181846 856
rect 182014 274 182490 856
rect 182658 274 183134 856
rect 183302 274 183778 856
rect 183946 274 184422 856
rect 184590 274 185066 856
rect 185234 274 185710 856
rect 185878 274 186354 856
rect 186522 274 186998 856
rect 187166 274 187642 856
rect 187810 274 188286 856
rect 188454 274 188930 856
rect 189098 274 189574 856
rect 189742 274 190218 856
rect 190386 274 190862 856
rect 191030 274 191506 856
rect 191674 274 192150 856
rect 192318 274 192794 856
rect 192962 274 193438 856
rect 193606 274 194082 856
rect 194250 274 194726 856
rect 194894 274 195370 856
rect 195538 274 196014 856
rect 196182 274 196658 856
rect 196826 274 197302 856
rect 197470 274 197946 856
rect 198114 274 198590 856
rect 198758 274 199234 856
rect 199402 274 199878 856
rect 200046 274 200522 856
rect 200690 274 201166 856
rect 201334 274 201810 856
rect 201978 274 202454 856
rect 202622 274 203098 856
rect 203266 274 203742 856
rect 203910 274 204386 856
rect 204554 274 205030 856
rect 205198 274 205674 856
rect 205842 274 206318 856
rect 206486 274 206962 856
rect 207130 274 207606 856
rect 207774 274 208250 856
rect 208418 274 208894 856
rect 209062 274 209538 856
rect 209706 274 210182 856
rect 210350 274 210826 856
rect 210994 274 211470 856
rect 211638 274 212114 856
rect 212282 274 212758 856
rect 212926 274 213402 856
rect 213570 274 214046 856
rect 214214 274 214690 856
rect 214858 274 215334 856
rect 215502 274 215978 856
rect 216146 274 216622 856
rect 216790 274 217266 856
rect 217434 274 217910 856
rect 218078 274 218554 856
rect 218722 274 219198 856
rect 219366 274 219842 856
rect 220010 274 220486 856
rect 220654 274 221130 856
rect 221298 274 221774 856
rect 221942 274 222418 856
rect 222586 274 223062 856
rect 223230 274 223706 856
rect 223874 274 224350 856
rect 224518 274 224994 856
rect 225162 274 225638 856
rect 225806 274 226282 856
rect 226450 274 226926 856
rect 227094 274 227570 856
rect 227738 274 228214 856
rect 228382 274 228858 856
rect 229026 274 229502 856
rect 229670 274 230146 856
rect 230314 274 230790 856
rect 230958 274 231434 856
rect 231602 274 232078 856
rect 232246 274 232722 856
rect 232890 274 233366 856
rect 233534 274 234010 856
rect 234178 274 234654 856
rect 234822 274 235298 856
rect 235466 274 235942 856
rect 236110 274 236586 856
rect 236754 274 237230 856
rect 237398 274 237874 856
rect 238042 274 238518 856
rect 238686 274 239162 856
rect 239330 274 239806 856
rect 239974 274 240450 856
rect 240618 274 241094 856
rect 241262 274 241738 856
rect 241906 274 242382 856
rect 242550 274 243026 856
rect 243194 274 243670 856
rect 243838 274 244314 856
rect 244482 274 244958 856
rect 245126 274 245602 856
rect 245770 274 246246 856
rect 246414 274 246890 856
rect 247058 274 247534 856
rect 247702 274 248178 856
rect 248346 274 248822 856
rect 248990 274 249466 856
rect 249634 274 250110 856
rect 250278 274 250754 856
rect 250922 274 251398 856
rect 251566 274 252042 856
rect 252210 274 252686 856
rect 252854 274 253330 856
rect 253498 274 253974 856
rect 254142 274 254618 856
rect 254786 274 255262 856
rect 255430 274 255906 856
rect 256074 274 256550 856
rect 256718 274 257194 856
rect 257362 274 257838 856
rect 258006 274 258482 856
rect 258650 274 259126 856
rect 259294 274 259770 856
rect 259938 274 260414 856
rect 260582 274 261058 856
rect 261226 274 261702 856
rect 261870 274 262346 856
rect 262514 274 262990 856
rect 263158 274 263634 856
rect 263802 274 264278 856
rect 264446 274 264922 856
rect 265090 274 265566 856
rect 265734 274 266210 856
rect 266378 274 266854 856
rect 267022 274 267498 856
rect 267666 274 268142 856
rect 268310 274 268786 856
rect 268954 274 269430 856
rect 269598 274 270074 856
rect 270242 274 270718 856
rect 270886 274 271362 856
rect 271530 274 272006 856
rect 272174 274 272650 856
rect 272818 274 273294 856
rect 273462 274 273938 856
rect 274106 274 274582 856
rect 274750 274 275226 856
rect 275394 274 275870 856
rect 276038 274 276514 856
rect 276682 274 277158 856
rect 277326 274 277802 856
rect 277970 274 278446 856
rect 278614 274 279090 856
rect 279258 274 279734 856
rect 279902 274 280378 856
rect 280546 274 281022 856
rect 281190 274 281666 856
rect 281834 274 282310 856
rect 282478 274 282954 856
rect 283122 274 283598 856
rect 283766 274 284242 856
rect 284410 274 284886 856
rect 285054 274 285530 856
rect 285698 274 286174 856
rect 286342 274 286818 856
rect 286986 274 287462 856
rect 287630 274 288106 856
rect 288274 274 288750 856
rect 288918 274 289394 856
rect 289562 274 290038 856
rect 290206 274 290682 856
rect 290850 274 291326 856
rect 291494 274 291970 856
rect 292138 274 292614 856
rect 292782 274 293258 856
rect 293426 274 293902 856
rect 294070 274 294546 856
rect 294714 274 295190 856
rect 295358 274 295834 856
rect 296002 274 296478 856
rect 296646 274 297122 856
rect 297290 274 297766 856
rect 297934 274 298410 856
rect 298578 274 299054 856
rect 299222 274 299698 856
rect 299866 274 300342 856
rect 300510 274 300986 856
rect 301154 274 301630 856
rect 301798 274 302274 856
rect 302442 274 302918 856
rect 303086 274 303562 856
rect 303730 274 304206 856
rect 304374 274 304850 856
rect 305018 274 305494 856
rect 305662 274 306138 856
rect 306306 274 306782 856
rect 306950 274 307426 856
rect 307594 274 308070 856
rect 308238 274 308714 856
rect 308882 274 309358 856
rect 309526 274 310002 856
rect 310170 274 310646 856
rect 310814 274 311290 856
rect 311458 274 311934 856
rect 312102 274 312578 856
rect 312746 274 313222 856
rect 313390 274 313866 856
rect 314034 274 314510 856
rect 314678 274 315154 856
rect 315322 274 315798 856
rect 315966 274 316442 856
rect 316610 274 317086 856
rect 317254 274 317730 856
rect 317898 274 318374 856
rect 318542 274 319018 856
rect 319186 274 319662 856
rect 319830 274 320306 856
rect 320474 274 320950 856
rect 321118 274 321594 856
rect 321762 274 322238 856
rect 322406 274 322882 856
rect 323050 274 323526 856
rect 323694 274 324170 856
rect 324338 274 324814 856
rect 324982 274 325458 856
rect 325626 274 326102 856
rect 326270 274 326746 856
rect 326914 274 327390 856
rect 327558 274 328034 856
rect 328202 274 328678 856
rect 328846 274 329322 856
rect 329490 274 329966 856
rect 330134 274 330610 856
rect 330778 274 331254 856
rect 331422 274 331898 856
rect 332066 274 332542 856
rect 332710 274 333186 856
rect 333354 274 333830 856
rect 333998 274 334474 856
rect 334642 274 335118 856
rect 335286 274 335762 856
rect 335930 274 336406 856
rect 336574 274 337050 856
rect 337218 274 337694 856
rect 337862 274 338338 856
rect 338506 274 358596 856
<< obsm3 >>
rect 381 444 357867 477665
<< metal4 >>
rect 4208 2128 4528 477680
rect 19568 2128 19888 477680
rect 34928 2128 35248 477680
rect 50288 2128 50608 477680
rect 65648 2128 65968 477680
rect 81008 2128 81328 477680
rect 96368 2128 96688 477680
rect 111728 2128 112048 477680
rect 127088 2128 127408 477680
rect 142448 2128 142768 477680
rect 157808 2128 158128 477680
rect 173168 2128 173488 477680
rect 188528 2128 188848 477680
rect 203888 2128 204208 477680
rect 219248 2128 219568 477680
rect 234608 2128 234928 477680
rect 249968 2128 250288 477680
rect 265328 2128 265648 477680
rect 280688 2128 281008 477680
rect 296048 2128 296368 477680
rect 311408 2128 311728 477680
rect 326768 2128 327088 477680
rect 342128 2128 342448 477680
rect 357488 2128 357808 477680
<< obsm4 >>
rect 427 2048 4128 476237
rect 4608 2048 19488 476237
rect 19968 2048 34848 476237
rect 35328 2048 50208 476237
rect 50688 2048 65568 476237
rect 66048 2048 80928 476237
rect 81408 2048 96288 476237
rect 96768 2048 111648 476237
rect 112128 2048 127008 476237
rect 127488 2048 142368 476237
rect 142848 2048 157728 476237
rect 158208 2048 173088 476237
rect 173568 2048 188448 476237
rect 188928 2048 203808 476237
rect 204288 2048 219168 476237
rect 219648 2048 234528 476237
rect 235008 2048 249888 476237
rect 250368 2048 265248 476237
rect 265728 2048 280608 476237
rect 281088 2048 295968 476237
rect 296448 2048 311328 476237
rect 311808 2048 326688 476237
rect 327168 2048 342048 476237
rect 342528 2048 348805 476237
rect 427 443 348805 2048
<< labels >>
rlabel metal2 s 3238 479200 3294 480000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 97078 479200 97134 480000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 106462 479200 106518 480000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 115846 479200 115902 480000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 125230 479200 125286 480000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 134614 479200 134670 480000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 143998 479200 144054 480000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 153382 479200 153438 480000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 162766 479200 162822 480000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 172150 479200 172206 480000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 181534 479200 181590 480000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12622 479200 12678 480000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 190918 479200 190974 480000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 200302 479200 200358 480000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 209686 479200 209742 480000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 219070 479200 219126 480000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 228454 479200 228510 480000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 237838 479200 237894 480000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 247222 479200 247278 480000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 256606 479200 256662 480000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 265990 479200 266046 480000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 275374 479200 275430 480000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22006 479200 22062 480000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 284758 479200 284814 480000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 294142 479200 294198 480000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 303526 479200 303582 480000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 312910 479200 312966 480000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 322294 479200 322350 480000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 331678 479200 331734 480000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 341062 479200 341118 480000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 350446 479200 350502 480000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 31390 479200 31446 480000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 40774 479200 40830 480000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 50158 479200 50214 480000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 59542 479200 59598 480000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 68926 479200 68982 480000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 78310 479200 78366 480000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 87694 479200 87750 480000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6366 479200 6422 480000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 100206 479200 100262 480000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 109590 479200 109646 480000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 118974 479200 119030 480000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 128358 479200 128414 480000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 137742 479200 137798 480000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 147126 479200 147182 480000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 156510 479200 156566 480000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 165894 479200 165950 480000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 175278 479200 175334 480000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 184662 479200 184718 480000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15750 479200 15806 480000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 194046 479200 194102 480000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 203430 479200 203486 480000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 212814 479200 212870 480000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 222198 479200 222254 480000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 231582 479200 231638 480000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 240966 479200 241022 480000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 250350 479200 250406 480000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 259734 479200 259790 480000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 269118 479200 269174 480000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 278502 479200 278558 480000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25134 479200 25190 480000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 287886 479200 287942 480000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 297270 479200 297326 480000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 306654 479200 306710 480000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 316038 479200 316094 480000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 325422 479200 325478 480000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 334806 479200 334862 480000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 344190 479200 344246 480000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 353574 479200 353630 480000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 34518 479200 34574 480000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 43902 479200 43958 480000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 53286 479200 53342 480000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 62670 479200 62726 480000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 72054 479200 72110 480000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 81438 479200 81494 480000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 90822 479200 90878 480000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9494 479200 9550 480000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 103334 479200 103390 480000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 112718 479200 112774 480000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 122102 479200 122158 480000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 131486 479200 131542 480000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 140870 479200 140926 480000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 150254 479200 150310 480000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 159638 479200 159694 480000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 169022 479200 169078 480000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 178406 479200 178462 480000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 187790 479200 187846 480000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 18878 479200 18934 480000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 197174 479200 197230 480000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 206558 479200 206614 480000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 215942 479200 215998 480000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 225326 479200 225382 480000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 234710 479200 234766 480000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 244094 479200 244150 480000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 253478 479200 253534 480000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 262862 479200 262918 480000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 272246 479200 272302 480000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 281630 479200 281686 480000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 28262 479200 28318 480000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 291014 479200 291070 480000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 300398 479200 300454 480000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 309782 479200 309838 480000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 319166 479200 319222 480000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 328550 479200 328606 480000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 337934 479200 337990 480000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 347318 479200 347374 480000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 356702 479200 356758 480000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 37646 479200 37702 480000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 47030 479200 47086 480000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 56414 479200 56470 480000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 65798 479200 65854 480000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 75182 479200 75238 480000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 84566 479200 84622 480000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 93950 479200 94006 480000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 337106 0 337162 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 337750 0 337806 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 338394 0 338450 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 288806 0 288862 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 290738 0 290794 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 296534 0 296590 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 298466 0 298522 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 302330 0 302386 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 304262 0 304318 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 308126 0 308182 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 310058 0 310114 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 311990 0 312046 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 313922 0 313978 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 317786 0 317842 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 319718 0 319774 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 323582 0 323638 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 325514 0 325570 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 327446 0 327502 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 333242 0 333298 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 335174 0 335230 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 263690 0 263746 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 271418 0 271474 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 275282 0 275338 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 279146 0 279202 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 285586 0 285642 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 287518 0 287574 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 289450 0 289506 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 291382 0 291438 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 293314 0 293370 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 295246 0 295302 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 297178 0 297234 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 299110 0 299166 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 302974 0 303030 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 306838 0 306894 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 308770 0 308826 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 310702 0 310758 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 312634 0 312690 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 314566 0 314622 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 316498 0 316554 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 320362 0 320418 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 324226 0 324282 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 326158 0 326214 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 328090 0 328146 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 331954 0 332010 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 333886 0 333942 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 335818 0 335874 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 185122 0 185178 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 192850 0 192906 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 194782 0 194838 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 204442 0 204498 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 206374 0 206430 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 208306 0 208362 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 210238 0 210294 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 212170 0 212226 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 216034 0 216090 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 217966 0 218022 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 225694 0 225750 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 227626 0 227682 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 233422 0 233478 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 235354 0 235410 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 237286 0 237342 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 241150 0 241206 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 245014 0 245070 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 246946 0 247002 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 250810 0 250866 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 258538 0 258594 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 270130 0 270186 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 272062 0 272118 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 273994 0 274050 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 275926 0 275982 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 279790 0 279846 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 286230 0 286286 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 290094 0 290150 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 292026 0 292082 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 295890 0 295946 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 305550 0 305606 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 307482 0 307538 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 309414 0 309470 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 311346 0 311402 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 313278 0 313334 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 317142 0 317198 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 319074 0 319130 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 321006 0 321062 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 326802 0 326858 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 328734 0 328790 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 330666 0 330722 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 234066 0 234122 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 235998 0 236054 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 243726 0 243782 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 264978 0 265034 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 266910 0 266966 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 268842 0 268898 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 270774 0 270830 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 282366 0 282422 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 477680 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 477680 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 21546 0 21602 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 360000 480000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 359065182
string GDS_FILE /home/htamas/progs/trainable-nn/openlane/trainable_nn/runs/22_09_12_18_06/results/signoff/trainable_nn.magic.gds
string GDS_START 1816374
<< end >>

