VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO trainable_nn
  CLASS BLOCK ;
  FOREIGN trainable_nn ;
  ORIGIN 0.000 0.000 ;
  SIZE 2200.000 BY 2800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 2796.000 34.410 2800.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 2796.000 600.210 2800.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 2796.000 656.790 2800.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 2796.000 713.370 2800.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 2796.000 769.950 2800.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 2796.000 826.530 2800.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 2796.000 883.110 2800.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 2796.000 939.690 2800.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 2796.000 996.270 2800.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 2796.000 1052.850 2800.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 2796.000 1109.430 2800.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 2796.000 90.990 2800.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 2796.000 1166.010 2800.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.310 2796.000 1222.590 2800.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 2796.000 1279.170 2800.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.470 2796.000 1335.750 2800.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.050 2796.000 1392.330 2800.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.630 2796.000 1448.910 2800.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.210 2796.000 1505.490 2800.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 2796.000 1562.070 2800.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 2796.000 1618.650 2800.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 2796.000 1675.230 2800.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 2796.000 147.570 2800.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 2796.000 1731.810 2800.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.110 2796.000 1788.390 2800.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.690 2796.000 1844.970 2800.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.270 2796.000 1901.550 2800.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 2796.000 1958.130 2800.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.430 2796.000 2014.710 2800.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.010 2796.000 2071.290 2800.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.590 2796.000 2127.870 2800.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 2796.000 204.150 2800.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 2796.000 260.730 2800.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 2796.000 317.310 2800.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 2796.000 373.890 2800.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 2796.000 430.470 2800.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 2796.000 487.050 2800.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 2796.000 543.630 2800.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 2796.000 53.270 2800.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 2796.000 619.070 2800.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 2796.000 675.650 2800.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 2796.000 732.230 2800.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 2796.000 788.810 2800.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 2796.000 845.390 2800.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 2796.000 901.970 2800.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 2796.000 958.550 2800.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 2796.000 1015.130 2800.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 2796.000 1071.710 2800.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 2796.000 1128.290 2800.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 2796.000 109.850 2800.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.590 2796.000 1184.870 2800.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 2796.000 1241.450 2800.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 2796.000 1298.030 2800.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.330 2796.000 1354.610 2800.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 2796.000 1411.190 2800.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.490 2796.000 1467.770 2800.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.070 2796.000 1524.350 2800.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 2796.000 1580.930 2800.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.230 2796.000 1637.510 2800.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 2796.000 1694.090 2800.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 2796.000 166.430 2800.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.390 2796.000 1750.670 2800.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.970 2796.000 1807.250 2800.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.550 2796.000 1863.830 2800.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.130 2796.000 1920.410 2800.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.710 2796.000 1976.990 2800.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.290 2796.000 2033.570 2800.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.870 2796.000 2090.150 2800.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.450 2796.000 2146.730 2800.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 2796.000 223.010 2800.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 2796.000 279.590 2800.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 2796.000 336.170 2800.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 2796.000 392.750 2800.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 2796.000 449.330 2800.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 2796.000 505.910 2800.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 2796.000 562.490 2800.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 2796.000 72.130 2800.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 2796.000 637.930 2800.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 2796.000 694.510 2800.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 2796.000 751.090 2800.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 2796.000 807.670 2800.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 2796.000 864.250 2800.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 2796.000 920.830 2800.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 2796.000 977.410 2800.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 2796.000 1033.990 2800.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 2796.000 1090.570 2800.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 2796.000 1147.150 2800.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 2796.000 128.710 2800.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 2796.000 1203.730 2800.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.030 2796.000 1260.310 2800.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.610 2796.000 1316.890 2800.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 2796.000 1373.470 2800.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 2796.000 1430.050 2800.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.350 2796.000 1486.630 2800.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 2796.000 1543.210 2800.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 2796.000 1599.790 2800.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 2796.000 1656.370 2800.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 2796.000 1712.950 2800.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 2796.000 185.290 2800.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.250 2796.000 1769.530 2800.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 2796.000 1826.110 2800.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.410 2796.000 1882.690 2800.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 2796.000 1939.270 2800.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.570 2796.000 1995.850 2800.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.150 2796.000 2052.430 2800.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.730 2796.000 2109.010 2800.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.310 2796.000 2165.590 2800.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 2796.000 241.870 2800.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 2796.000 298.450 2800.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 2796.000 355.030 2800.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 2796.000 411.610 2800.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 2796.000 468.190 2800.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 2796.000 524.770 2800.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 2796.000 581.350 2800.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2110.110 0.000 2110.390 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.250 0.000 2114.530 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.390 0.000 2118.670 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.350 0.000 1762.630 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.770 0.000 1775.050 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.610 0.000 1799.890 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.030 0.000 1812.310 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.450 0.000 1824.730 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.870 0.000 1837.150 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 0.000 1849.570 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 0.000 1861.990 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.550 0.000 1886.830 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.970 0.000 1899.250 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.390 0.000 1911.670 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.810 0.000 1924.090 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.230 0.000 1936.510 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.650 0.000 1948.930 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 0.000 1986.190 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.330 0.000 1998.610 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.750 0.000 2011.030 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.170 0.000 2023.450 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.590 0.000 2035.870 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 0.000 2048.290 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 0.000 2060.710 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.850 0.000 2073.130 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.270 0.000 2085.550 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.690 0.000 2097.970 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 0.000 868.390 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 0.000 1042.270 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 0.000 1154.050 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 0.000 1203.730 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 0.000 1216.150 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 0.000 1228.570 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 0.000 1240.990 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 0.000 1290.670 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 0.000 1303.090 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.230 0.000 1315.510 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 0.000 1327.930 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 0.000 1340.350 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.910 0.000 1365.190 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.330 0.000 1377.610 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 0.000 1390.030 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.170 0.000 1402.450 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 0.000 1427.290 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 0.000 1452.130 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 0.000 1464.550 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.790 0.000 1539.070 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 0.000 1588.750 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 0.000 1626.010 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.150 0.000 1638.430 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 0.000 1663.270 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 0.000 1688.110 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 0.000 1712.950 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 0.000 1725.370 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.930 0.000 1750.210 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.490 0.000 1766.770 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.910 0.000 1779.190 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.750 0.000 1804.030 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.590 0.000 1828.870 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.010 0.000 1841.290 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 0.000 1853.710 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.850 0.000 1866.130 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.270 0.000 1878.550 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 0.000 1890.970 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 0.000 1903.390 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.950 0.000 1928.230 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.370 0.000 1940.650 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.790 0.000 1953.070 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.210 0.000 1965.490 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.630 0.000 1977.910 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.470 0.000 2002.750 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.890 0.000 2015.170 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.310 0.000 2027.590 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.730 0.000 2040.010 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.570 0.000 2064.850 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.410 0.000 2089.690 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.830 0.000 2102.110 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 0.000 959.470 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 0.000 1083.670 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 0.000 1158.190 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 0.000 1170.610 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 0.000 1245.130 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 0.000 1282.390 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 0.000 1307.230 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 0.000 1369.330 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.150 0.000 1431.430 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 0.000 1443.850 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.830 0.000 1481.110 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.250 0.000 1493.530 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.670 0.000 1505.950 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 0.000 1518.370 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 0.000 1530.790 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 0.000 1592.890 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 0.000 1617.730 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.870 0.000 1630.150 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 0.000 1654.990 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 0.000 1667.410 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550 0.000 1679.830 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 0.000 1704.670 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 0.000 1754.350 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 0.000 1770.910 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 0.000 1783.330 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.470 0.000 1795.750 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.310 0.000 1820.590 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.730 0.000 1833.010 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.990 0.000 1870.270 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.410 0.000 1882.690 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.250 0.000 1907.530 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 0.000 1919.950 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.510 0.000 1944.790 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.930 0.000 1957.210 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.770 0.000 1982.050 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.190 0.000 1994.470 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.610 0.000 2006.890 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.450 0.000 2031.730 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.870 0.000 2044.150 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2056.290 0.000 2056.570 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.710 0.000 2068.990 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.130 0.000 2081.410 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.550 0.000 2093.830 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 0.000 826.990 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 0.000 1025.710 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 0.000 1162.330 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 0.000 1261.690 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 0.000 1286.530 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 0.000 1298.950 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 0.000 1311.370 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 0.000 1385.890 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 0.000 1398.310 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 0.000 1460.410 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 0.000 1472.830 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 0.000 1485.250 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.810 0.000 1510.090 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.230 0.000 1522.510 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 0.000 1534.930 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.070 0.000 1547.350 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 0.000 1559.770 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 0.000 1572.190 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 0.000 1597.030 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 0.000 1609.450 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 0.000 1621.870 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.010 0.000 1634.290 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.430 0.000 1646.710 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 0.000 1659.130 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 0.000 1683.970 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.110 0.000 1696.390 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 0.000 1708.810 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.950 0.000 1721.230 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.370 0.000 1733.650 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 0.000 1746.070 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2788.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2788.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2788.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 2786.585 2194.390 2788.190 ;
        RECT 5.330 2781.145 2194.390 2783.975 ;
        RECT 5.330 2775.705 2194.390 2778.535 ;
        RECT 5.330 2770.265 2194.390 2773.095 ;
        RECT 5.330 2764.825 2194.390 2767.655 ;
        RECT 5.330 2759.385 2194.390 2762.215 ;
        RECT 5.330 2753.945 2194.390 2756.775 ;
        RECT 5.330 2748.505 2194.390 2751.335 ;
        RECT 5.330 2743.065 2194.390 2745.895 ;
        RECT 5.330 2737.625 2194.390 2740.455 ;
        RECT 5.330 2732.185 2194.390 2735.015 ;
        RECT 5.330 2726.745 2194.390 2729.575 ;
        RECT 5.330 2721.305 2194.390 2724.135 ;
        RECT 5.330 2715.865 2194.390 2718.695 ;
        RECT 5.330 2710.425 2194.390 2713.255 ;
        RECT 5.330 2704.985 2194.390 2707.815 ;
        RECT 5.330 2699.545 2194.390 2702.375 ;
        RECT 5.330 2694.105 2194.390 2696.935 ;
        RECT 5.330 2688.665 2194.390 2691.495 ;
        RECT 5.330 2683.225 2194.390 2686.055 ;
        RECT 5.330 2677.785 2194.390 2680.615 ;
        RECT 5.330 2672.345 2194.390 2675.175 ;
        RECT 5.330 2666.905 2194.390 2669.735 ;
        RECT 5.330 2661.465 2194.390 2664.295 ;
        RECT 5.330 2656.025 2194.390 2658.855 ;
        RECT 5.330 2650.585 2194.390 2653.415 ;
        RECT 5.330 2645.145 2194.390 2647.975 ;
        RECT 5.330 2639.705 2194.390 2642.535 ;
        RECT 5.330 2634.265 2194.390 2637.095 ;
        RECT 5.330 2628.825 2194.390 2631.655 ;
        RECT 5.330 2623.385 2194.390 2626.215 ;
        RECT 5.330 2617.945 2194.390 2620.775 ;
        RECT 5.330 2612.505 2194.390 2615.335 ;
        RECT 5.330 2607.065 2194.390 2609.895 ;
        RECT 5.330 2601.625 2194.390 2604.455 ;
        RECT 5.330 2596.185 2194.390 2599.015 ;
        RECT 5.330 2590.745 2194.390 2593.575 ;
        RECT 5.330 2585.305 2194.390 2588.135 ;
        RECT 5.330 2579.865 2194.390 2582.695 ;
        RECT 5.330 2574.425 2194.390 2577.255 ;
        RECT 5.330 2568.985 2194.390 2571.815 ;
        RECT 5.330 2563.545 2194.390 2566.375 ;
        RECT 5.330 2558.105 2194.390 2560.935 ;
        RECT 5.330 2552.665 2194.390 2555.495 ;
        RECT 5.330 2547.225 2194.390 2550.055 ;
        RECT 5.330 2541.785 2194.390 2544.615 ;
        RECT 5.330 2536.345 2194.390 2539.175 ;
        RECT 5.330 2530.905 2194.390 2533.735 ;
        RECT 5.330 2525.465 2194.390 2528.295 ;
        RECT 5.330 2520.025 2194.390 2522.855 ;
        RECT 5.330 2514.585 2194.390 2517.415 ;
        RECT 5.330 2509.145 2194.390 2511.975 ;
        RECT 5.330 2503.705 2194.390 2506.535 ;
        RECT 5.330 2498.265 2194.390 2501.095 ;
        RECT 5.330 2492.825 2194.390 2495.655 ;
        RECT 5.330 2487.385 2194.390 2490.215 ;
        RECT 5.330 2481.945 2194.390 2484.775 ;
        RECT 5.330 2476.505 2194.390 2479.335 ;
        RECT 5.330 2471.065 2194.390 2473.895 ;
        RECT 5.330 2465.625 2194.390 2468.455 ;
        RECT 5.330 2460.185 2194.390 2463.015 ;
        RECT 5.330 2454.745 2194.390 2457.575 ;
        RECT 5.330 2449.305 2194.390 2452.135 ;
        RECT 5.330 2443.865 2194.390 2446.695 ;
        RECT 5.330 2438.425 2194.390 2441.255 ;
        RECT 5.330 2432.985 2194.390 2435.815 ;
        RECT 5.330 2427.545 2194.390 2430.375 ;
        RECT 5.330 2422.105 2194.390 2424.935 ;
        RECT 5.330 2416.665 2194.390 2419.495 ;
        RECT 5.330 2411.225 2194.390 2414.055 ;
        RECT 5.330 2405.785 2194.390 2408.615 ;
        RECT 5.330 2400.345 2194.390 2403.175 ;
        RECT 5.330 2394.905 2194.390 2397.735 ;
        RECT 5.330 2389.465 2194.390 2392.295 ;
        RECT 5.330 2384.025 2194.390 2386.855 ;
        RECT 5.330 2378.585 2194.390 2381.415 ;
        RECT 5.330 2373.145 2194.390 2375.975 ;
        RECT 5.330 2367.705 2194.390 2370.535 ;
        RECT 5.330 2362.265 2194.390 2365.095 ;
        RECT 5.330 2356.825 2194.390 2359.655 ;
        RECT 5.330 2351.385 2194.390 2354.215 ;
        RECT 5.330 2345.945 2194.390 2348.775 ;
        RECT 5.330 2340.505 2194.390 2343.335 ;
        RECT 5.330 2335.065 2194.390 2337.895 ;
        RECT 5.330 2329.625 2194.390 2332.455 ;
        RECT 5.330 2324.185 2194.390 2327.015 ;
        RECT 5.330 2318.745 2194.390 2321.575 ;
        RECT 5.330 2313.305 2194.390 2316.135 ;
        RECT 5.330 2307.865 2194.390 2310.695 ;
        RECT 5.330 2302.425 2194.390 2305.255 ;
        RECT 5.330 2296.985 2194.390 2299.815 ;
        RECT 5.330 2291.545 2194.390 2294.375 ;
        RECT 5.330 2286.105 2194.390 2288.935 ;
        RECT 5.330 2280.665 2194.390 2283.495 ;
        RECT 5.330 2275.225 2194.390 2278.055 ;
        RECT 5.330 2269.785 2194.390 2272.615 ;
        RECT 5.330 2264.345 2194.390 2267.175 ;
        RECT 5.330 2258.905 2194.390 2261.735 ;
        RECT 5.330 2253.465 2194.390 2256.295 ;
        RECT 5.330 2248.025 2194.390 2250.855 ;
        RECT 5.330 2242.585 2194.390 2245.415 ;
        RECT 5.330 2237.145 2194.390 2239.975 ;
        RECT 5.330 2231.705 2194.390 2234.535 ;
        RECT 5.330 2226.265 2194.390 2229.095 ;
        RECT 5.330 2220.825 2194.390 2223.655 ;
        RECT 5.330 2215.385 2194.390 2218.215 ;
        RECT 5.330 2209.945 2194.390 2212.775 ;
        RECT 5.330 2204.505 2194.390 2207.335 ;
        RECT 5.330 2199.065 2194.390 2201.895 ;
        RECT 5.330 2193.625 2194.390 2196.455 ;
        RECT 5.330 2188.185 2194.390 2191.015 ;
        RECT 5.330 2182.745 2194.390 2185.575 ;
        RECT 5.330 2177.305 2194.390 2180.135 ;
        RECT 5.330 2171.865 2194.390 2174.695 ;
        RECT 5.330 2166.425 2194.390 2169.255 ;
        RECT 5.330 2160.985 2194.390 2163.815 ;
        RECT 5.330 2155.545 2194.390 2158.375 ;
        RECT 5.330 2150.105 2194.390 2152.935 ;
        RECT 5.330 2144.665 2194.390 2147.495 ;
        RECT 5.330 2139.225 2194.390 2142.055 ;
        RECT 5.330 2133.785 2194.390 2136.615 ;
        RECT 5.330 2128.345 2194.390 2131.175 ;
        RECT 5.330 2122.905 2194.390 2125.735 ;
        RECT 5.330 2117.465 2194.390 2120.295 ;
        RECT 5.330 2112.025 2194.390 2114.855 ;
        RECT 5.330 2106.585 2194.390 2109.415 ;
        RECT 5.330 2101.145 2194.390 2103.975 ;
        RECT 5.330 2095.705 2194.390 2098.535 ;
        RECT 5.330 2090.265 2194.390 2093.095 ;
        RECT 5.330 2084.825 2194.390 2087.655 ;
        RECT 5.330 2079.385 2194.390 2082.215 ;
        RECT 5.330 2073.945 2194.390 2076.775 ;
        RECT 5.330 2068.505 2194.390 2071.335 ;
        RECT 5.330 2063.065 2194.390 2065.895 ;
        RECT 5.330 2057.625 2194.390 2060.455 ;
        RECT 5.330 2052.185 2194.390 2055.015 ;
        RECT 5.330 2046.745 2194.390 2049.575 ;
        RECT 5.330 2041.305 2194.390 2044.135 ;
        RECT 5.330 2035.865 2194.390 2038.695 ;
        RECT 5.330 2030.425 2194.390 2033.255 ;
        RECT 5.330 2024.985 2194.390 2027.815 ;
        RECT 5.330 2019.545 2194.390 2022.375 ;
        RECT 5.330 2014.105 2194.390 2016.935 ;
        RECT 5.330 2008.665 2194.390 2011.495 ;
        RECT 5.330 2003.225 2194.390 2006.055 ;
        RECT 5.330 1997.785 2194.390 2000.615 ;
        RECT 5.330 1992.345 2194.390 1995.175 ;
        RECT 5.330 1986.905 2194.390 1989.735 ;
        RECT 5.330 1981.465 2194.390 1984.295 ;
        RECT 5.330 1976.025 2194.390 1978.855 ;
        RECT 5.330 1970.585 2194.390 1973.415 ;
        RECT 5.330 1965.145 2194.390 1967.975 ;
        RECT 5.330 1959.705 2194.390 1962.535 ;
        RECT 5.330 1954.265 2194.390 1957.095 ;
        RECT 5.330 1948.825 2194.390 1951.655 ;
        RECT 5.330 1943.385 2194.390 1946.215 ;
        RECT 5.330 1937.945 2194.390 1940.775 ;
        RECT 5.330 1932.505 2194.390 1935.335 ;
        RECT 5.330 1927.065 2194.390 1929.895 ;
        RECT 5.330 1921.625 2194.390 1924.455 ;
        RECT 5.330 1916.185 2194.390 1919.015 ;
        RECT 5.330 1910.745 2194.390 1913.575 ;
        RECT 5.330 1905.305 2194.390 1908.135 ;
        RECT 5.330 1899.865 2194.390 1902.695 ;
        RECT 5.330 1894.425 2194.390 1897.255 ;
        RECT 5.330 1888.985 2194.390 1891.815 ;
        RECT 5.330 1883.545 2194.390 1886.375 ;
        RECT 5.330 1878.105 2194.390 1880.935 ;
        RECT 5.330 1872.665 2194.390 1875.495 ;
        RECT 5.330 1867.225 2194.390 1870.055 ;
        RECT 5.330 1861.785 2194.390 1864.615 ;
        RECT 5.330 1856.345 2194.390 1859.175 ;
        RECT 5.330 1850.905 2194.390 1853.735 ;
        RECT 5.330 1845.465 2194.390 1848.295 ;
        RECT 5.330 1840.025 2194.390 1842.855 ;
        RECT 5.330 1834.585 2194.390 1837.415 ;
        RECT 5.330 1829.145 2194.390 1831.975 ;
        RECT 5.330 1823.705 2194.390 1826.535 ;
        RECT 5.330 1818.265 2194.390 1821.095 ;
        RECT 5.330 1812.825 2194.390 1815.655 ;
        RECT 5.330 1807.385 2194.390 1810.215 ;
        RECT 5.330 1801.945 2194.390 1804.775 ;
        RECT 5.330 1796.505 2194.390 1799.335 ;
        RECT 5.330 1791.065 2194.390 1793.895 ;
        RECT 5.330 1785.625 2194.390 1788.455 ;
        RECT 5.330 1780.185 2194.390 1783.015 ;
        RECT 5.330 1774.745 2194.390 1777.575 ;
        RECT 5.330 1769.305 2194.390 1772.135 ;
        RECT 5.330 1763.865 2194.390 1766.695 ;
        RECT 5.330 1758.425 2194.390 1761.255 ;
        RECT 5.330 1752.985 2194.390 1755.815 ;
        RECT 5.330 1747.545 2194.390 1750.375 ;
        RECT 5.330 1742.105 2194.390 1744.935 ;
        RECT 5.330 1736.665 2194.390 1739.495 ;
        RECT 5.330 1731.225 2194.390 1734.055 ;
        RECT 5.330 1725.785 2194.390 1728.615 ;
        RECT 5.330 1720.345 2194.390 1723.175 ;
        RECT 5.330 1714.905 2194.390 1717.735 ;
        RECT 5.330 1709.465 2194.390 1712.295 ;
        RECT 5.330 1704.025 2194.390 1706.855 ;
        RECT 5.330 1698.585 2194.390 1701.415 ;
        RECT 5.330 1693.145 2194.390 1695.975 ;
        RECT 5.330 1687.705 2194.390 1690.535 ;
        RECT 5.330 1682.265 2194.390 1685.095 ;
        RECT 5.330 1676.825 2194.390 1679.655 ;
        RECT 5.330 1671.385 2194.390 1674.215 ;
        RECT 5.330 1665.945 2194.390 1668.775 ;
        RECT 5.330 1660.505 2194.390 1663.335 ;
        RECT 5.330 1655.065 2194.390 1657.895 ;
        RECT 5.330 1649.625 2194.390 1652.455 ;
        RECT 5.330 1644.185 2194.390 1647.015 ;
        RECT 5.330 1638.745 2194.390 1641.575 ;
        RECT 5.330 1633.305 2194.390 1636.135 ;
        RECT 5.330 1627.865 2194.390 1630.695 ;
        RECT 5.330 1622.425 2194.390 1625.255 ;
        RECT 5.330 1616.985 2194.390 1619.815 ;
        RECT 5.330 1611.545 2194.390 1614.375 ;
        RECT 5.330 1606.105 2194.390 1608.935 ;
        RECT 5.330 1600.665 2194.390 1603.495 ;
        RECT 5.330 1595.225 2194.390 1598.055 ;
        RECT 5.330 1589.785 2194.390 1592.615 ;
        RECT 5.330 1584.345 2194.390 1587.175 ;
        RECT 5.330 1578.905 2194.390 1581.735 ;
        RECT 5.330 1573.465 2194.390 1576.295 ;
        RECT 5.330 1568.025 2194.390 1570.855 ;
        RECT 5.330 1562.585 2194.390 1565.415 ;
        RECT 5.330 1557.145 2194.390 1559.975 ;
        RECT 5.330 1551.705 2194.390 1554.535 ;
        RECT 5.330 1546.265 2194.390 1549.095 ;
        RECT 5.330 1540.825 2194.390 1543.655 ;
        RECT 5.330 1535.385 2194.390 1538.215 ;
        RECT 5.330 1529.945 2194.390 1532.775 ;
        RECT 5.330 1524.505 2194.390 1527.335 ;
        RECT 5.330 1519.065 2194.390 1521.895 ;
        RECT 5.330 1513.625 2194.390 1516.455 ;
        RECT 5.330 1508.185 2194.390 1511.015 ;
        RECT 5.330 1502.745 2194.390 1505.575 ;
        RECT 5.330 1497.305 2194.390 1500.135 ;
        RECT 5.330 1491.865 2194.390 1494.695 ;
        RECT 5.330 1486.425 2194.390 1489.255 ;
        RECT 5.330 1480.985 2194.390 1483.815 ;
        RECT 5.330 1475.545 2194.390 1478.375 ;
        RECT 5.330 1470.105 2194.390 1472.935 ;
        RECT 5.330 1464.665 2194.390 1467.495 ;
        RECT 5.330 1459.225 2194.390 1462.055 ;
        RECT 5.330 1453.785 2194.390 1456.615 ;
        RECT 5.330 1448.345 2194.390 1451.175 ;
        RECT 5.330 1442.905 2194.390 1445.735 ;
        RECT 5.330 1437.465 2194.390 1440.295 ;
        RECT 5.330 1432.025 2194.390 1434.855 ;
        RECT 5.330 1426.585 2194.390 1429.415 ;
        RECT 5.330 1421.145 2194.390 1423.975 ;
        RECT 5.330 1415.705 2194.390 1418.535 ;
        RECT 5.330 1410.265 2194.390 1413.095 ;
        RECT 5.330 1404.825 2194.390 1407.655 ;
        RECT 5.330 1399.385 2194.390 1402.215 ;
        RECT 5.330 1393.945 2194.390 1396.775 ;
        RECT 5.330 1388.505 2194.390 1391.335 ;
        RECT 5.330 1383.065 2194.390 1385.895 ;
        RECT 5.330 1377.625 2194.390 1380.455 ;
        RECT 5.330 1372.185 2194.390 1375.015 ;
        RECT 5.330 1366.745 2194.390 1369.575 ;
        RECT 5.330 1361.305 2194.390 1364.135 ;
        RECT 5.330 1355.865 2194.390 1358.695 ;
        RECT 5.330 1350.425 2194.390 1353.255 ;
        RECT 5.330 1344.985 2194.390 1347.815 ;
        RECT 5.330 1339.545 2194.390 1342.375 ;
        RECT 5.330 1334.105 2194.390 1336.935 ;
        RECT 5.330 1328.665 2194.390 1331.495 ;
        RECT 5.330 1323.225 2194.390 1326.055 ;
        RECT 5.330 1317.785 2194.390 1320.615 ;
        RECT 5.330 1312.345 2194.390 1315.175 ;
        RECT 5.330 1306.905 2194.390 1309.735 ;
        RECT 5.330 1301.465 2194.390 1304.295 ;
        RECT 5.330 1296.025 2194.390 1298.855 ;
        RECT 5.330 1290.585 2194.390 1293.415 ;
        RECT 5.330 1285.145 2194.390 1287.975 ;
        RECT 5.330 1279.705 2194.390 1282.535 ;
        RECT 5.330 1274.265 2194.390 1277.095 ;
        RECT 5.330 1268.825 2194.390 1271.655 ;
        RECT 5.330 1263.385 2194.390 1266.215 ;
        RECT 5.330 1257.945 2194.390 1260.775 ;
        RECT 5.330 1252.505 2194.390 1255.335 ;
        RECT 5.330 1247.065 2194.390 1249.895 ;
        RECT 5.330 1241.625 2194.390 1244.455 ;
        RECT 5.330 1236.185 2194.390 1239.015 ;
        RECT 5.330 1230.745 2194.390 1233.575 ;
        RECT 5.330 1225.305 2194.390 1228.135 ;
        RECT 5.330 1219.865 2194.390 1222.695 ;
        RECT 5.330 1214.425 2194.390 1217.255 ;
        RECT 5.330 1208.985 2194.390 1211.815 ;
        RECT 5.330 1203.545 2194.390 1206.375 ;
        RECT 5.330 1198.105 2194.390 1200.935 ;
        RECT 5.330 1192.665 2194.390 1195.495 ;
        RECT 5.330 1187.225 2194.390 1190.055 ;
        RECT 5.330 1181.785 2194.390 1184.615 ;
        RECT 5.330 1176.345 2194.390 1179.175 ;
        RECT 5.330 1170.905 2194.390 1173.735 ;
        RECT 5.330 1165.465 2194.390 1168.295 ;
        RECT 5.330 1160.025 2194.390 1162.855 ;
        RECT 5.330 1154.585 2194.390 1157.415 ;
        RECT 5.330 1149.145 2194.390 1151.975 ;
        RECT 5.330 1143.705 2194.390 1146.535 ;
        RECT 5.330 1138.265 2194.390 1141.095 ;
        RECT 5.330 1132.825 2194.390 1135.655 ;
        RECT 5.330 1127.385 2194.390 1130.215 ;
        RECT 5.330 1121.945 2194.390 1124.775 ;
        RECT 5.330 1116.505 2194.390 1119.335 ;
        RECT 5.330 1111.065 2194.390 1113.895 ;
        RECT 5.330 1105.625 2194.390 1108.455 ;
        RECT 5.330 1100.185 2194.390 1103.015 ;
        RECT 5.330 1094.745 2194.390 1097.575 ;
        RECT 5.330 1089.305 2194.390 1092.135 ;
        RECT 5.330 1083.865 2194.390 1086.695 ;
        RECT 5.330 1078.425 2194.390 1081.255 ;
        RECT 5.330 1072.985 2194.390 1075.815 ;
        RECT 5.330 1067.545 2194.390 1070.375 ;
        RECT 5.330 1062.105 2194.390 1064.935 ;
        RECT 5.330 1056.665 2194.390 1059.495 ;
        RECT 5.330 1051.225 2194.390 1054.055 ;
        RECT 5.330 1045.785 2194.390 1048.615 ;
        RECT 5.330 1040.345 2194.390 1043.175 ;
        RECT 5.330 1034.905 2194.390 1037.735 ;
        RECT 5.330 1029.465 2194.390 1032.295 ;
        RECT 5.330 1024.025 2194.390 1026.855 ;
        RECT 5.330 1018.585 2194.390 1021.415 ;
        RECT 5.330 1013.145 2194.390 1015.975 ;
        RECT 5.330 1007.705 2194.390 1010.535 ;
        RECT 5.330 1002.265 2194.390 1005.095 ;
        RECT 5.330 996.825 2194.390 999.655 ;
        RECT 5.330 991.385 2194.390 994.215 ;
        RECT 5.330 985.945 2194.390 988.775 ;
        RECT 5.330 980.505 2194.390 983.335 ;
        RECT 5.330 975.065 2194.390 977.895 ;
        RECT 5.330 969.625 2194.390 972.455 ;
        RECT 5.330 964.185 2194.390 967.015 ;
        RECT 5.330 958.745 2194.390 961.575 ;
        RECT 5.330 953.305 2194.390 956.135 ;
        RECT 5.330 947.865 2194.390 950.695 ;
        RECT 5.330 942.425 2194.390 945.255 ;
        RECT 5.330 936.985 2194.390 939.815 ;
        RECT 5.330 931.545 2194.390 934.375 ;
        RECT 5.330 926.105 2194.390 928.935 ;
        RECT 5.330 920.665 2194.390 923.495 ;
        RECT 5.330 915.225 2194.390 918.055 ;
        RECT 5.330 909.785 2194.390 912.615 ;
        RECT 5.330 904.345 2194.390 907.175 ;
        RECT 5.330 898.905 2194.390 901.735 ;
        RECT 5.330 893.465 2194.390 896.295 ;
        RECT 5.330 888.025 2194.390 890.855 ;
        RECT 5.330 882.585 2194.390 885.415 ;
        RECT 5.330 877.145 2194.390 879.975 ;
        RECT 5.330 871.705 2194.390 874.535 ;
        RECT 5.330 866.265 2194.390 869.095 ;
        RECT 5.330 860.825 2194.390 863.655 ;
        RECT 5.330 855.385 2194.390 858.215 ;
        RECT 5.330 849.945 2194.390 852.775 ;
        RECT 5.330 844.505 2194.390 847.335 ;
        RECT 5.330 839.065 2194.390 841.895 ;
        RECT 5.330 833.625 2194.390 836.455 ;
        RECT 5.330 828.185 2194.390 831.015 ;
        RECT 5.330 822.745 2194.390 825.575 ;
        RECT 5.330 817.305 2194.390 820.135 ;
        RECT 5.330 811.865 2194.390 814.695 ;
        RECT 5.330 806.425 2194.390 809.255 ;
        RECT 5.330 800.985 2194.390 803.815 ;
        RECT 5.330 795.545 2194.390 798.375 ;
        RECT 5.330 790.105 2194.390 792.935 ;
        RECT 5.330 784.665 2194.390 787.495 ;
        RECT 5.330 779.225 2194.390 782.055 ;
        RECT 5.330 773.785 2194.390 776.615 ;
        RECT 5.330 768.345 2194.390 771.175 ;
        RECT 5.330 762.905 2194.390 765.735 ;
        RECT 5.330 757.465 2194.390 760.295 ;
        RECT 5.330 752.025 2194.390 754.855 ;
        RECT 5.330 746.585 2194.390 749.415 ;
        RECT 5.330 741.145 2194.390 743.975 ;
        RECT 5.330 735.705 2194.390 738.535 ;
        RECT 5.330 730.265 2194.390 733.095 ;
        RECT 5.330 724.825 2194.390 727.655 ;
        RECT 5.330 719.385 2194.390 722.215 ;
        RECT 5.330 713.945 2194.390 716.775 ;
        RECT 5.330 708.505 2194.390 711.335 ;
        RECT 5.330 703.065 2194.390 705.895 ;
        RECT 5.330 697.625 2194.390 700.455 ;
        RECT 5.330 692.185 2194.390 695.015 ;
        RECT 5.330 686.745 2194.390 689.575 ;
        RECT 5.330 681.305 2194.390 684.135 ;
        RECT 5.330 675.865 2194.390 678.695 ;
        RECT 5.330 670.425 2194.390 673.255 ;
        RECT 5.330 664.985 2194.390 667.815 ;
        RECT 5.330 659.545 2194.390 662.375 ;
        RECT 5.330 654.105 2194.390 656.935 ;
        RECT 5.330 648.665 2194.390 651.495 ;
        RECT 5.330 643.225 2194.390 646.055 ;
        RECT 5.330 637.785 2194.390 640.615 ;
        RECT 5.330 632.345 2194.390 635.175 ;
        RECT 5.330 626.905 2194.390 629.735 ;
        RECT 5.330 621.465 2194.390 624.295 ;
        RECT 5.330 616.025 2194.390 618.855 ;
        RECT 5.330 610.585 2194.390 613.415 ;
        RECT 5.330 605.145 2194.390 607.975 ;
        RECT 5.330 599.705 2194.390 602.535 ;
        RECT 5.330 594.265 2194.390 597.095 ;
        RECT 5.330 588.825 2194.390 591.655 ;
        RECT 5.330 583.385 2194.390 586.215 ;
        RECT 5.330 577.945 2194.390 580.775 ;
        RECT 5.330 572.505 2194.390 575.335 ;
        RECT 5.330 567.065 2194.390 569.895 ;
        RECT 5.330 561.625 2194.390 564.455 ;
        RECT 5.330 556.185 2194.390 559.015 ;
        RECT 5.330 550.745 2194.390 553.575 ;
        RECT 5.330 545.305 2194.390 548.135 ;
        RECT 5.330 539.865 2194.390 542.695 ;
        RECT 5.330 534.425 2194.390 537.255 ;
        RECT 5.330 528.985 2194.390 531.815 ;
        RECT 5.330 523.545 2194.390 526.375 ;
        RECT 5.330 518.105 2194.390 520.935 ;
        RECT 5.330 512.665 2194.390 515.495 ;
        RECT 5.330 507.225 2194.390 510.055 ;
        RECT 5.330 501.785 2194.390 504.615 ;
        RECT 5.330 496.345 2194.390 499.175 ;
        RECT 5.330 490.905 2194.390 493.735 ;
        RECT 5.330 485.465 2194.390 488.295 ;
        RECT 5.330 480.025 2194.390 482.855 ;
        RECT 5.330 474.585 2194.390 477.415 ;
        RECT 5.330 469.145 2194.390 471.975 ;
        RECT 5.330 463.705 2194.390 466.535 ;
        RECT 5.330 458.265 2194.390 461.095 ;
        RECT 5.330 452.825 2194.390 455.655 ;
        RECT 5.330 447.385 2194.390 450.215 ;
        RECT 5.330 441.945 2194.390 444.775 ;
        RECT 5.330 436.505 2194.390 439.335 ;
        RECT 5.330 431.065 2194.390 433.895 ;
        RECT 5.330 425.625 2194.390 428.455 ;
        RECT 5.330 420.185 2194.390 423.015 ;
        RECT 5.330 414.745 2194.390 417.575 ;
        RECT 5.330 409.305 2194.390 412.135 ;
        RECT 5.330 403.865 2194.390 406.695 ;
        RECT 5.330 398.425 2194.390 401.255 ;
        RECT 5.330 392.985 2194.390 395.815 ;
        RECT 5.330 387.545 2194.390 390.375 ;
        RECT 5.330 382.105 2194.390 384.935 ;
        RECT 5.330 376.665 2194.390 379.495 ;
        RECT 5.330 371.225 2194.390 374.055 ;
        RECT 5.330 365.785 2194.390 368.615 ;
        RECT 5.330 360.345 2194.390 363.175 ;
        RECT 5.330 354.905 2194.390 357.735 ;
        RECT 5.330 349.465 2194.390 352.295 ;
        RECT 5.330 344.025 2194.390 346.855 ;
        RECT 5.330 338.585 2194.390 341.415 ;
        RECT 5.330 333.145 2194.390 335.975 ;
        RECT 5.330 327.705 2194.390 330.535 ;
        RECT 5.330 322.265 2194.390 325.095 ;
        RECT 5.330 316.825 2194.390 319.655 ;
        RECT 5.330 311.385 2194.390 314.215 ;
        RECT 5.330 305.945 2194.390 308.775 ;
        RECT 5.330 300.505 2194.390 303.335 ;
        RECT 5.330 295.065 2194.390 297.895 ;
        RECT 5.330 289.625 2194.390 292.455 ;
        RECT 5.330 284.185 2194.390 287.015 ;
        RECT 5.330 278.745 2194.390 281.575 ;
        RECT 5.330 273.305 2194.390 276.135 ;
        RECT 5.330 267.865 2194.390 270.695 ;
        RECT 5.330 262.425 2194.390 265.255 ;
        RECT 5.330 256.985 2194.390 259.815 ;
        RECT 5.330 251.545 2194.390 254.375 ;
        RECT 5.330 246.105 2194.390 248.935 ;
        RECT 5.330 240.665 2194.390 243.495 ;
        RECT 5.330 235.225 2194.390 238.055 ;
        RECT 5.330 229.785 2194.390 232.615 ;
        RECT 5.330 224.345 2194.390 227.175 ;
        RECT 5.330 218.905 2194.390 221.735 ;
        RECT 5.330 213.465 2194.390 216.295 ;
        RECT 5.330 208.025 2194.390 210.855 ;
        RECT 5.330 202.585 2194.390 205.415 ;
        RECT 5.330 197.145 2194.390 199.975 ;
        RECT 5.330 191.705 2194.390 194.535 ;
        RECT 5.330 186.265 2194.390 189.095 ;
        RECT 5.330 180.825 2194.390 183.655 ;
        RECT 5.330 175.385 2194.390 178.215 ;
        RECT 5.330 169.945 2194.390 172.775 ;
        RECT 5.330 164.505 2194.390 167.335 ;
        RECT 5.330 159.065 2194.390 161.895 ;
        RECT 5.330 153.625 2194.390 156.455 ;
        RECT 5.330 148.185 2194.390 151.015 ;
        RECT 5.330 142.745 2194.390 145.575 ;
        RECT 5.330 137.305 2194.390 140.135 ;
        RECT 5.330 131.865 2194.390 134.695 ;
        RECT 5.330 126.425 2194.390 129.255 ;
        RECT 5.330 120.985 2194.390 123.815 ;
        RECT 5.330 115.545 2194.390 118.375 ;
        RECT 5.330 110.105 2194.390 112.935 ;
        RECT 5.330 104.665 2194.390 107.495 ;
        RECT 5.330 99.225 2194.390 102.055 ;
        RECT 5.330 93.785 2194.390 96.615 ;
        RECT 5.330 88.345 2194.390 91.175 ;
        RECT 5.330 82.905 2194.390 85.735 ;
        RECT 5.330 77.465 2194.390 80.295 ;
        RECT 5.330 72.025 2194.390 74.855 ;
        RECT 5.330 66.585 2194.390 69.415 ;
        RECT 5.330 61.145 2194.390 63.975 ;
        RECT 5.330 55.705 2194.390 58.535 ;
        RECT 5.330 50.265 2194.390 53.095 ;
        RECT 5.330 44.825 2194.390 47.655 ;
        RECT 5.330 39.385 2194.390 42.215 ;
        RECT 5.330 33.945 2194.390 36.775 ;
        RECT 5.330 28.505 2194.390 31.335 ;
        RECT 5.330 23.065 2194.390 25.895 ;
        RECT 5.330 17.625 2194.390 20.455 ;
        RECT 5.330 12.185 2194.390 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 2194.200 2788.085 ;
      LAYER met1 ;
        RECT 5.520 0.720 2195.050 2788.240 ;
      LAYER met2 ;
        RECT 7.000 2795.720 33.850 2796.570 ;
        RECT 34.690 2795.720 52.710 2796.570 ;
        RECT 53.550 2795.720 71.570 2796.570 ;
        RECT 72.410 2795.720 90.430 2796.570 ;
        RECT 91.270 2795.720 109.290 2796.570 ;
        RECT 110.130 2795.720 128.150 2796.570 ;
        RECT 128.990 2795.720 147.010 2796.570 ;
        RECT 147.850 2795.720 165.870 2796.570 ;
        RECT 166.710 2795.720 184.730 2796.570 ;
        RECT 185.570 2795.720 203.590 2796.570 ;
        RECT 204.430 2795.720 222.450 2796.570 ;
        RECT 223.290 2795.720 241.310 2796.570 ;
        RECT 242.150 2795.720 260.170 2796.570 ;
        RECT 261.010 2795.720 279.030 2796.570 ;
        RECT 279.870 2795.720 297.890 2796.570 ;
        RECT 298.730 2795.720 316.750 2796.570 ;
        RECT 317.590 2795.720 335.610 2796.570 ;
        RECT 336.450 2795.720 354.470 2796.570 ;
        RECT 355.310 2795.720 373.330 2796.570 ;
        RECT 374.170 2795.720 392.190 2796.570 ;
        RECT 393.030 2795.720 411.050 2796.570 ;
        RECT 411.890 2795.720 429.910 2796.570 ;
        RECT 430.750 2795.720 448.770 2796.570 ;
        RECT 449.610 2795.720 467.630 2796.570 ;
        RECT 468.470 2795.720 486.490 2796.570 ;
        RECT 487.330 2795.720 505.350 2796.570 ;
        RECT 506.190 2795.720 524.210 2796.570 ;
        RECT 525.050 2795.720 543.070 2796.570 ;
        RECT 543.910 2795.720 561.930 2796.570 ;
        RECT 562.770 2795.720 580.790 2796.570 ;
        RECT 581.630 2795.720 599.650 2796.570 ;
        RECT 600.490 2795.720 618.510 2796.570 ;
        RECT 619.350 2795.720 637.370 2796.570 ;
        RECT 638.210 2795.720 656.230 2796.570 ;
        RECT 657.070 2795.720 675.090 2796.570 ;
        RECT 675.930 2795.720 693.950 2796.570 ;
        RECT 694.790 2795.720 712.810 2796.570 ;
        RECT 713.650 2795.720 731.670 2796.570 ;
        RECT 732.510 2795.720 750.530 2796.570 ;
        RECT 751.370 2795.720 769.390 2796.570 ;
        RECT 770.230 2795.720 788.250 2796.570 ;
        RECT 789.090 2795.720 807.110 2796.570 ;
        RECT 807.950 2795.720 825.970 2796.570 ;
        RECT 826.810 2795.720 844.830 2796.570 ;
        RECT 845.670 2795.720 863.690 2796.570 ;
        RECT 864.530 2795.720 882.550 2796.570 ;
        RECT 883.390 2795.720 901.410 2796.570 ;
        RECT 902.250 2795.720 920.270 2796.570 ;
        RECT 921.110 2795.720 939.130 2796.570 ;
        RECT 939.970 2795.720 957.990 2796.570 ;
        RECT 958.830 2795.720 976.850 2796.570 ;
        RECT 977.690 2795.720 995.710 2796.570 ;
        RECT 996.550 2795.720 1014.570 2796.570 ;
        RECT 1015.410 2795.720 1033.430 2796.570 ;
        RECT 1034.270 2795.720 1052.290 2796.570 ;
        RECT 1053.130 2795.720 1071.150 2796.570 ;
        RECT 1071.990 2795.720 1090.010 2796.570 ;
        RECT 1090.850 2795.720 1108.870 2796.570 ;
        RECT 1109.710 2795.720 1127.730 2796.570 ;
        RECT 1128.570 2795.720 1146.590 2796.570 ;
        RECT 1147.430 2795.720 1165.450 2796.570 ;
        RECT 1166.290 2795.720 1184.310 2796.570 ;
        RECT 1185.150 2795.720 1203.170 2796.570 ;
        RECT 1204.010 2795.720 1222.030 2796.570 ;
        RECT 1222.870 2795.720 1240.890 2796.570 ;
        RECT 1241.730 2795.720 1259.750 2796.570 ;
        RECT 1260.590 2795.720 1278.610 2796.570 ;
        RECT 1279.450 2795.720 1297.470 2796.570 ;
        RECT 1298.310 2795.720 1316.330 2796.570 ;
        RECT 1317.170 2795.720 1335.190 2796.570 ;
        RECT 1336.030 2795.720 1354.050 2796.570 ;
        RECT 1354.890 2795.720 1372.910 2796.570 ;
        RECT 1373.750 2795.720 1391.770 2796.570 ;
        RECT 1392.610 2795.720 1410.630 2796.570 ;
        RECT 1411.470 2795.720 1429.490 2796.570 ;
        RECT 1430.330 2795.720 1448.350 2796.570 ;
        RECT 1449.190 2795.720 1467.210 2796.570 ;
        RECT 1468.050 2795.720 1486.070 2796.570 ;
        RECT 1486.910 2795.720 1504.930 2796.570 ;
        RECT 1505.770 2795.720 1523.790 2796.570 ;
        RECT 1524.630 2795.720 1542.650 2796.570 ;
        RECT 1543.490 2795.720 1561.510 2796.570 ;
        RECT 1562.350 2795.720 1580.370 2796.570 ;
        RECT 1581.210 2795.720 1599.230 2796.570 ;
        RECT 1600.070 2795.720 1618.090 2796.570 ;
        RECT 1618.930 2795.720 1636.950 2796.570 ;
        RECT 1637.790 2795.720 1655.810 2796.570 ;
        RECT 1656.650 2795.720 1674.670 2796.570 ;
        RECT 1675.510 2795.720 1693.530 2796.570 ;
        RECT 1694.370 2795.720 1712.390 2796.570 ;
        RECT 1713.230 2795.720 1731.250 2796.570 ;
        RECT 1732.090 2795.720 1750.110 2796.570 ;
        RECT 1750.950 2795.720 1768.970 2796.570 ;
        RECT 1769.810 2795.720 1787.830 2796.570 ;
        RECT 1788.670 2795.720 1806.690 2796.570 ;
        RECT 1807.530 2795.720 1825.550 2796.570 ;
        RECT 1826.390 2795.720 1844.410 2796.570 ;
        RECT 1845.250 2795.720 1863.270 2796.570 ;
        RECT 1864.110 2795.720 1882.130 2796.570 ;
        RECT 1882.970 2795.720 1900.990 2796.570 ;
        RECT 1901.830 2795.720 1919.850 2796.570 ;
        RECT 1920.690 2795.720 1938.710 2796.570 ;
        RECT 1939.550 2795.720 1957.570 2796.570 ;
        RECT 1958.410 2795.720 1976.430 2796.570 ;
        RECT 1977.270 2795.720 1995.290 2796.570 ;
        RECT 1996.130 2795.720 2014.150 2796.570 ;
        RECT 2014.990 2795.720 2033.010 2796.570 ;
        RECT 2033.850 2795.720 2051.870 2796.570 ;
        RECT 2052.710 2795.720 2070.730 2796.570 ;
        RECT 2071.570 2795.720 2089.590 2796.570 ;
        RECT 2090.430 2795.720 2108.450 2796.570 ;
        RECT 2109.290 2795.720 2127.310 2796.570 ;
        RECT 2128.150 2795.720 2146.170 2796.570 ;
        RECT 2147.010 2795.720 2165.030 2796.570 ;
        RECT 2165.870 2795.720 2195.030 2796.570 ;
        RECT 7.000 4.280 2195.030 2795.720 ;
        RECT 7.000 0.690 81.230 4.280 ;
        RECT 82.070 0.690 85.370 4.280 ;
        RECT 86.210 0.690 89.510 4.280 ;
        RECT 90.350 0.690 93.650 4.280 ;
        RECT 94.490 0.690 97.790 4.280 ;
        RECT 98.630 0.690 101.930 4.280 ;
        RECT 102.770 0.690 106.070 4.280 ;
        RECT 106.910 0.690 110.210 4.280 ;
        RECT 111.050 0.690 114.350 4.280 ;
        RECT 115.190 0.690 118.490 4.280 ;
        RECT 119.330 0.690 122.630 4.280 ;
        RECT 123.470 0.690 126.770 4.280 ;
        RECT 127.610 0.690 130.910 4.280 ;
        RECT 131.750 0.690 135.050 4.280 ;
        RECT 135.890 0.690 139.190 4.280 ;
        RECT 140.030 0.690 143.330 4.280 ;
        RECT 144.170 0.690 147.470 4.280 ;
        RECT 148.310 0.690 151.610 4.280 ;
        RECT 152.450 0.690 155.750 4.280 ;
        RECT 156.590 0.690 159.890 4.280 ;
        RECT 160.730 0.690 164.030 4.280 ;
        RECT 164.870 0.690 168.170 4.280 ;
        RECT 169.010 0.690 172.310 4.280 ;
        RECT 173.150 0.690 176.450 4.280 ;
        RECT 177.290 0.690 180.590 4.280 ;
        RECT 181.430 0.690 184.730 4.280 ;
        RECT 185.570 0.690 188.870 4.280 ;
        RECT 189.710 0.690 193.010 4.280 ;
        RECT 193.850 0.690 197.150 4.280 ;
        RECT 197.990 0.690 201.290 4.280 ;
        RECT 202.130 0.690 205.430 4.280 ;
        RECT 206.270 0.690 209.570 4.280 ;
        RECT 210.410 0.690 213.710 4.280 ;
        RECT 214.550 0.690 217.850 4.280 ;
        RECT 218.690 0.690 221.990 4.280 ;
        RECT 222.830 0.690 226.130 4.280 ;
        RECT 226.970 0.690 230.270 4.280 ;
        RECT 231.110 0.690 234.410 4.280 ;
        RECT 235.250 0.690 238.550 4.280 ;
        RECT 239.390 0.690 242.690 4.280 ;
        RECT 243.530 0.690 246.830 4.280 ;
        RECT 247.670 0.690 250.970 4.280 ;
        RECT 251.810 0.690 255.110 4.280 ;
        RECT 255.950 0.690 259.250 4.280 ;
        RECT 260.090 0.690 263.390 4.280 ;
        RECT 264.230 0.690 267.530 4.280 ;
        RECT 268.370 0.690 271.670 4.280 ;
        RECT 272.510 0.690 275.810 4.280 ;
        RECT 276.650 0.690 279.950 4.280 ;
        RECT 280.790 0.690 284.090 4.280 ;
        RECT 284.930 0.690 288.230 4.280 ;
        RECT 289.070 0.690 292.370 4.280 ;
        RECT 293.210 0.690 296.510 4.280 ;
        RECT 297.350 0.690 300.650 4.280 ;
        RECT 301.490 0.690 304.790 4.280 ;
        RECT 305.630 0.690 308.930 4.280 ;
        RECT 309.770 0.690 313.070 4.280 ;
        RECT 313.910 0.690 317.210 4.280 ;
        RECT 318.050 0.690 321.350 4.280 ;
        RECT 322.190 0.690 325.490 4.280 ;
        RECT 326.330 0.690 329.630 4.280 ;
        RECT 330.470 0.690 333.770 4.280 ;
        RECT 334.610 0.690 337.910 4.280 ;
        RECT 338.750 0.690 342.050 4.280 ;
        RECT 342.890 0.690 346.190 4.280 ;
        RECT 347.030 0.690 350.330 4.280 ;
        RECT 351.170 0.690 354.470 4.280 ;
        RECT 355.310 0.690 358.610 4.280 ;
        RECT 359.450 0.690 362.750 4.280 ;
        RECT 363.590 0.690 366.890 4.280 ;
        RECT 367.730 0.690 371.030 4.280 ;
        RECT 371.870 0.690 375.170 4.280 ;
        RECT 376.010 0.690 379.310 4.280 ;
        RECT 380.150 0.690 383.450 4.280 ;
        RECT 384.290 0.690 387.590 4.280 ;
        RECT 388.430 0.690 391.730 4.280 ;
        RECT 392.570 0.690 395.870 4.280 ;
        RECT 396.710 0.690 400.010 4.280 ;
        RECT 400.850 0.690 404.150 4.280 ;
        RECT 404.990 0.690 408.290 4.280 ;
        RECT 409.130 0.690 412.430 4.280 ;
        RECT 413.270 0.690 416.570 4.280 ;
        RECT 417.410 0.690 420.710 4.280 ;
        RECT 421.550 0.690 424.850 4.280 ;
        RECT 425.690 0.690 428.990 4.280 ;
        RECT 429.830 0.690 433.130 4.280 ;
        RECT 433.970 0.690 437.270 4.280 ;
        RECT 438.110 0.690 441.410 4.280 ;
        RECT 442.250 0.690 445.550 4.280 ;
        RECT 446.390 0.690 449.690 4.280 ;
        RECT 450.530 0.690 453.830 4.280 ;
        RECT 454.670 0.690 457.970 4.280 ;
        RECT 458.810 0.690 462.110 4.280 ;
        RECT 462.950 0.690 466.250 4.280 ;
        RECT 467.090 0.690 470.390 4.280 ;
        RECT 471.230 0.690 474.530 4.280 ;
        RECT 475.370 0.690 478.670 4.280 ;
        RECT 479.510 0.690 482.810 4.280 ;
        RECT 483.650 0.690 486.950 4.280 ;
        RECT 487.790 0.690 491.090 4.280 ;
        RECT 491.930 0.690 495.230 4.280 ;
        RECT 496.070 0.690 499.370 4.280 ;
        RECT 500.210 0.690 503.510 4.280 ;
        RECT 504.350 0.690 507.650 4.280 ;
        RECT 508.490 0.690 511.790 4.280 ;
        RECT 512.630 0.690 515.930 4.280 ;
        RECT 516.770 0.690 520.070 4.280 ;
        RECT 520.910 0.690 524.210 4.280 ;
        RECT 525.050 0.690 528.350 4.280 ;
        RECT 529.190 0.690 532.490 4.280 ;
        RECT 533.330 0.690 536.630 4.280 ;
        RECT 537.470 0.690 540.770 4.280 ;
        RECT 541.610 0.690 544.910 4.280 ;
        RECT 545.750 0.690 549.050 4.280 ;
        RECT 549.890 0.690 553.190 4.280 ;
        RECT 554.030 0.690 557.330 4.280 ;
        RECT 558.170 0.690 561.470 4.280 ;
        RECT 562.310 0.690 565.610 4.280 ;
        RECT 566.450 0.690 569.750 4.280 ;
        RECT 570.590 0.690 573.890 4.280 ;
        RECT 574.730 0.690 578.030 4.280 ;
        RECT 578.870 0.690 582.170 4.280 ;
        RECT 583.010 0.690 586.310 4.280 ;
        RECT 587.150 0.690 590.450 4.280 ;
        RECT 591.290 0.690 594.590 4.280 ;
        RECT 595.430 0.690 598.730 4.280 ;
        RECT 599.570 0.690 602.870 4.280 ;
        RECT 603.710 0.690 607.010 4.280 ;
        RECT 607.850 0.690 611.150 4.280 ;
        RECT 611.990 0.690 615.290 4.280 ;
        RECT 616.130 0.690 619.430 4.280 ;
        RECT 620.270 0.690 623.570 4.280 ;
        RECT 624.410 0.690 627.710 4.280 ;
        RECT 628.550 0.690 631.850 4.280 ;
        RECT 632.690 0.690 635.990 4.280 ;
        RECT 636.830 0.690 640.130 4.280 ;
        RECT 640.970 0.690 644.270 4.280 ;
        RECT 645.110 0.690 648.410 4.280 ;
        RECT 649.250 0.690 652.550 4.280 ;
        RECT 653.390 0.690 656.690 4.280 ;
        RECT 657.530 0.690 660.830 4.280 ;
        RECT 661.670 0.690 664.970 4.280 ;
        RECT 665.810 0.690 669.110 4.280 ;
        RECT 669.950 0.690 673.250 4.280 ;
        RECT 674.090 0.690 677.390 4.280 ;
        RECT 678.230 0.690 681.530 4.280 ;
        RECT 682.370 0.690 685.670 4.280 ;
        RECT 686.510 0.690 689.810 4.280 ;
        RECT 690.650 0.690 693.950 4.280 ;
        RECT 694.790 0.690 698.090 4.280 ;
        RECT 698.930 0.690 702.230 4.280 ;
        RECT 703.070 0.690 706.370 4.280 ;
        RECT 707.210 0.690 710.510 4.280 ;
        RECT 711.350 0.690 714.650 4.280 ;
        RECT 715.490 0.690 718.790 4.280 ;
        RECT 719.630 0.690 722.930 4.280 ;
        RECT 723.770 0.690 727.070 4.280 ;
        RECT 727.910 0.690 731.210 4.280 ;
        RECT 732.050 0.690 735.350 4.280 ;
        RECT 736.190 0.690 739.490 4.280 ;
        RECT 740.330 0.690 743.630 4.280 ;
        RECT 744.470 0.690 747.770 4.280 ;
        RECT 748.610 0.690 751.910 4.280 ;
        RECT 752.750 0.690 756.050 4.280 ;
        RECT 756.890 0.690 760.190 4.280 ;
        RECT 761.030 0.690 764.330 4.280 ;
        RECT 765.170 0.690 768.470 4.280 ;
        RECT 769.310 0.690 772.610 4.280 ;
        RECT 773.450 0.690 776.750 4.280 ;
        RECT 777.590 0.690 780.890 4.280 ;
        RECT 781.730 0.690 785.030 4.280 ;
        RECT 785.870 0.690 789.170 4.280 ;
        RECT 790.010 0.690 793.310 4.280 ;
        RECT 794.150 0.690 797.450 4.280 ;
        RECT 798.290 0.690 801.590 4.280 ;
        RECT 802.430 0.690 805.730 4.280 ;
        RECT 806.570 0.690 809.870 4.280 ;
        RECT 810.710 0.690 814.010 4.280 ;
        RECT 814.850 0.690 818.150 4.280 ;
        RECT 818.990 0.690 822.290 4.280 ;
        RECT 823.130 0.690 826.430 4.280 ;
        RECT 827.270 0.690 830.570 4.280 ;
        RECT 831.410 0.690 834.710 4.280 ;
        RECT 835.550 0.690 838.850 4.280 ;
        RECT 839.690 0.690 842.990 4.280 ;
        RECT 843.830 0.690 847.130 4.280 ;
        RECT 847.970 0.690 851.270 4.280 ;
        RECT 852.110 0.690 855.410 4.280 ;
        RECT 856.250 0.690 859.550 4.280 ;
        RECT 860.390 0.690 863.690 4.280 ;
        RECT 864.530 0.690 867.830 4.280 ;
        RECT 868.670 0.690 871.970 4.280 ;
        RECT 872.810 0.690 876.110 4.280 ;
        RECT 876.950 0.690 880.250 4.280 ;
        RECT 881.090 0.690 884.390 4.280 ;
        RECT 885.230 0.690 888.530 4.280 ;
        RECT 889.370 0.690 892.670 4.280 ;
        RECT 893.510 0.690 896.810 4.280 ;
        RECT 897.650 0.690 900.950 4.280 ;
        RECT 901.790 0.690 905.090 4.280 ;
        RECT 905.930 0.690 909.230 4.280 ;
        RECT 910.070 0.690 913.370 4.280 ;
        RECT 914.210 0.690 917.510 4.280 ;
        RECT 918.350 0.690 921.650 4.280 ;
        RECT 922.490 0.690 925.790 4.280 ;
        RECT 926.630 0.690 929.930 4.280 ;
        RECT 930.770 0.690 934.070 4.280 ;
        RECT 934.910 0.690 938.210 4.280 ;
        RECT 939.050 0.690 942.350 4.280 ;
        RECT 943.190 0.690 946.490 4.280 ;
        RECT 947.330 0.690 950.630 4.280 ;
        RECT 951.470 0.690 954.770 4.280 ;
        RECT 955.610 0.690 958.910 4.280 ;
        RECT 959.750 0.690 963.050 4.280 ;
        RECT 963.890 0.690 967.190 4.280 ;
        RECT 968.030 0.690 971.330 4.280 ;
        RECT 972.170 0.690 975.470 4.280 ;
        RECT 976.310 0.690 979.610 4.280 ;
        RECT 980.450 0.690 983.750 4.280 ;
        RECT 984.590 0.690 987.890 4.280 ;
        RECT 988.730 0.690 992.030 4.280 ;
        RECT 992.870 0.690 996.170 4.280 ;
        RECT 997.010 0.690 1000.310 4.280 ;
        RECT 1001.150 0.690 1004.450 4.280 ;
        RECT 1005.290 0.690 1008.590 4.280 ;
        RECT 1009.430 0.690 1012.730 4.280 ;
        RECT 1013.570 0.690 1016.870 4.280 ;
        RECT 1017.710 0.690 1021.010 4.280 ;
        RECT 1021.850 0.690 1025.150 4.280 ;
        RECT 1025.990 0.690 1029.290 4.280 ;
        RECT 1030.130 0.690 1033.430 4.280 ;
        RECT 1034.270 0.690 1037.570 4.280 ;
        RECT 1038.410 0.690 1041.710 4.280 ;
        RECT 1042.550 0.690 1045.850 4.280 ;
        RECT 1046.690 0.690 1049.990 4.280 ;
        RECT 1050.830 0.690 1054.130 4.280 ;
        RECT 1054.970 0.690 1058.270 4.280 ;
        RECT 1059.110 0.690 1062.410 4.280 ;
        RECT 1063.250 0.690 1066.550 4.280 ;
        RECT 1067.390 0.690 1070.690 4.280 ;
        RECT 1071.530 0.690 1074.830 4.280 ;
        RECT 1075.670 0.690 1078.970 4.280 ;
        RECT 1079.810 0.690 1083.110 4.280 ;
        RECT 1083.950 0.690 1087.250 4.280 ;
        RECT 1088.090 0.690 1091.390 4.280 ;
        RECT 1092.230 0.690 1095.530 4.280 ;
        RECT 1096.370 0.690 1099.670 4.280 ;
        RECT 1100.510 0.690 1103.810 4.280 ;
        RECT 1104.650 0.690 1107.950 4.280 ;
        RECT 1108.790 0.690 1112.090 4.280 ;
        RECT 1112.930 0.690 1116.230 4.280 ;
        RECT 1117.070 0.690 1120.370 4.280 ;
        RECT 1121.210 0.690 1124.510 4.280 ;
        RECT 1125.350 0.690 1128.650 4.280 ;
        RECT 1129.490 0.690 1132.790 4.280 ;
        RECT 1133.630 0.690 1136.930 4.280 ;
        RECT 1137.770 0.690 1141.070 4.280 ;
        RECT 1141.910 0.690 1145.210 4.280 ;
        RECT 1146.050 0.690 1149.350 4.280 ;
        RECT 1150.190 0.690 1153.490 4.280 ;
        RECT 1154.330 0.690 1157.630 4.280 ;
        RECT 1158.470 0.690 1161.770 4.280 ;
        RECT 1162.610 0.690 1165.910 4.280 ;
        RECT 1166.750 0.690 1170.050 4.280 ;
        RECT 1170.890 0.690 1174.190 4.280 ;
        RECT 1175.030 0.690 1178.330 4.280 ;
        RECT 1179.170 0.690 1182.470 4.280 ;
        RECT 1183.310 0.690 1186.610 4.280 ;
        RECT 1187.450 0.690 1190.750 4.280 ;
        RECT 1191.590 0.690 1194.890 4.280 ;
        RECT 1195.730 0.690 1199.030 4.280 ;
        RECT 1199.870 0.690 1203.170 4.280 ;
        RECT 1204.010 0.690 1207.310 4.280 ;
        RECT 1208.150 0.690 1211.450 4.280 ;
        RECT 1212.290 0.690 1215.590 4.280 ;
        RECT 1216.430 0.690 1219.730 4.280 ;
        RECT 1220.570 0.690 1223.870 4.280 ;
        RECT 1224.710 0.690 1228.010 4.280 ;
        RECT 1228.850 0.690 1232.150 4.280 ;
        RECT 1232.990 0.690 1236.290 4.280 ;
        RECT 1237.130 0.690 1240.430 4.280 ;
        RECT 1241.270 0.690 1244.570 4.280 ;
        RECT 1245.410 0.690 1248.710 4.280 ;
        RECT 1249.550 0.690 1252.850 4.280 ;
        RECT 1253.690 0.690 1256.990 4.280 ;
        RECT 1257.830 0.690 1261.130 4.280 ;
        RECT 1261.970 0.690 1265.270 4.280 ;
        RECT 1266.110 0.690 1269.410 4.280 ;
        RECT 1270.250 0.690 1273.550 4.280 ;
        RECT 1274.390 0.690 1277.690 4.280 ;
        RECT 1278.530 0.690 1281.830 4.280 ;
        RECT 1282.670 0.690 1285.970 4.280 ;
        RECT 1286.810 0.690 1290.110 4.280 ;
        RECT 1290.950 0.690 1294.250 4.280 ;
        RECT 1295.090 0.690 1298.390 4.280 ;
        RECT 1299.230 0.690 1302.530 4.280 ;
        RECT 1303.370 0.690 1306.670 4.280 ;
        RECT 1307.510 0.690 1310.810 4.280 ;
        RECT 1311.650 0.690 1314.950 4.280 ;
        RECT 1315.790 0.690 1319.090 4.280 ;
        RECT 1319.930 0.690 1323.230 4.280 ;
        RECT 1324.070 0.690 1327.370 4.280 ;
        RECT 1328.210 0.690 1331.510 4.280 ;
        RECT 1332.350 0.690 1335.650 4.280 ;
        RECT 1336.490 0.690 1339.790 4.280 ;
        RECT 1340.630 0.690 1343.930 4.280 ;
        RECT 1344.770 0.690 1348.070 4.280 ;
        RECT 1348.910 0.690 1352.210 4.280 ;
        RECT 1353.050 0.690 1356.350 4.280 ;
        RECT 1357.190 0.690 1360.490 4.280 ;
        RECT 1361.330 0.690 1364.630 4.280 ;
        RECT 1365.470 0.690 1368.770 4.280 ;
        RECT 1369.610 0.690 1372.910 4.280 ;
        RECT 1373.750 0.690 1377.050 4.280 ;
        RECT 1377.890 0.690 1381.190 4.280 ;
        RECT 1382.030 0.690 1385.330 4.280 ;
        RECT 1386.170 0.690 1389.470 4.280 ;
        RECT 1390.310 0.690 1393.610 4.280 ;
        RECT 1394.450 0.690 1397.750 4.280 ;
        RECT 1398.590 0.690 1401.890 4.280 ;
        RECT 1402.730 0.690 1406.030 4.280 ;
        RECT 1406.870 0.690 1410.170 4.280 ;
        RECT 1411.010 0.690 1414.310 4.280 ;
        RECT 1415.150 0.690 1418.450 4.280 ;
        RECT 1419.290 0.690 1422.590 4.280 ;
        RECT 1423.430 0.690 1426.730 4.280 ;
        RECT 1427.570 0.690 1430.870 4.280 ;
        RECT 1431.710 0.690 1435.010 4.280 ;
        RECT 1435.850 0.690 1439.150 4.280 ;
        RECT 1439.990 0.690 1443.290 4.280 ;
        RECT 1444.130 0.690 1447.430 4.280 ;
        RECT 1448.270 0.690 1451.570 4.280 ;
        RECT 1452.410 0.690 1455.710 4.280 ;
        RECT 1456.550 0.690 1459.850 4.280 ;
        RECT 1460.690 0.690 1463.990 4.280 ;
        RECT 1464.830 0.690 1468.130 4.280 ;
        RECT 1468.970 0.690 1472.270 4.280 ;
        RECT 1473.110 0.690 1476.410 4.280 ;
        RECT 1477.250 0.690 1480.550 4.280 ;
        RECT 1481.390 0.690 1484.690 4.280 ;
        RECT 1485.530 0.690 1488.830 4.280 ;
        RECT 1489.670 0.690 1492.970 4.280 ;
        RECT 1493.810 0.690 1497.110 4.280 ;
        RECT 1497.950 0.690 1501.250 4.280 ;
        RECT 1502.090 0.690 1505.390 4.280 ;
        RECT 1506.230 0.690 1509.530 4.280 ;
        RECT 1510.370 0.690 1513.670 4.280 ;
        RECT 1514.510 0.690 1517.810 4.280 ;
        RECT 1518.650 0.690 1521.950 4.280 ;
        RECT 1522.790 0.690 1526.090 4.280 ;
        RECT 1526.930 0.690 1530.230 4.280 ;
        RECT 1531.070 0.690 1534.370 4.280 ;
        RECT 1535.210 0.690 1538.510 4.280 ;
        RECT 1539.350 0.690 1542.650 4.280 ;
        RECT 1543.490 0.690 1546.790 4.280 ;
        RECT 1547.630 0.690 1550.930 4.280 ;
        RECT 1551.770 0.690 1555.070 4.280 ;
        RECT 1555.910 0.690 1559.210 4.280 ;
        RECT 1560.050 0.690 1563.350 4.280 ;
        RECT 1564.190 0.690 1567.490 4.280 ;
        RECT 1568.330 0.690 1571.630 4.280 ;
        RECT 1572.470 0.690 1575.770 4.280 ;
        RECT 1576.610 0.690 1579.910 4.280 ;
        RECT 1580.750 0.690 1584.050 4.280 ;
        RECT 1584.890 0.690 1588.190 4.280 ;
        RECT 1589.030 0.690 1592.330 4.280 ;
        RECT 1593.170 0.690 1596.470 4.280 ;
        RECT 1597.310 0.690 1600.610 4.280 ;
        RECT 1601.450 0.690 1604.750 4.280 ;
        RECT 1605.590 0.690 1608.890 4.280 ;
        RECT 1609.730 0.690 1613.030 4.280 ;
        RECT 1613.870 0.690 1617.170 4.280 ;
        RECT 1618.010 0.690 1621.310 4.280 ;
        RECT 1622.150 0.690 1625.450 4.280 ;
        RECT 1626.290 0.690 1629.590 4.280 ;
        RECT 1630.430 0.690 1633.730 4.280 ;
        RECT 1634.570 0.690 1637.870 4.280 ;
        RECT 1638.710 0.690 1642.010 4.280 ;
        RECT 1642.850 0.690 1646.150 4.280 ;
        RECT 1646.990 0.690 1650.290 4.280 ;
        RECT 1651.130 0.690 1654.430 4.280 ;
        RECT 1655.270 0.690 1658.570 4.280 ;
        RECT 1659.410 0.690 1662.710 4.280 ;
        RECT 1663.550 0.690 1666.850 4.280 ;
        RECT 1667.690 0.690 1670.990 4.280 ;
        RECT 1671.830 0.690 1675.130 4.280 ;
        RECT 1675.970 0.690 1679.270 4.280 ;
        RECT 1680.110 0.690 1683.410 4.280 ;
        RECT 1684.250 0.690 1687.550 4.280 ;
        RECT 1688.390 0.690 1691.690 4.280 ;
        RECT 1692.530 0.690 1695.830 4.280 ;
        RECT 1696.670 0.690 1699.970 4.280 ;
        RECT 1700.810 0.690 1704.110 4.280 ;
        RECT 1704.950 0.690 1708.250 4.280 ;
        RECT 1709.090 0.690 1712.390 4.280 ;
        RECT 1713.230 0.690 1716.530 4.280 ;
        RECT 1717.370 0.690 1720.670 4.280 ;
        RECT 1721.510 0.690 1724.810 4.280 ;
        RECT 1725.650 0.690 1728.950 4.280 ;
        RECT 1729.790 0.690 1733.090 4.280 ;
        RECT 1733.930 0.690 1737.230 4.280 ;
        RECT 1738.070 0.690 1741.370 4.280 ;
        RECT 1742.210 0.690 1745.510 4.280 ;
        RECT 1746.350 0.690 1749.650 4.280 ;
        RECT 1750.490 0.690 1753.790 4.280 ;
        RECT 1754.630 0.690 1757.930 4.280 ;
        RECT 1758.770 0.690 1762.070 4.280 ;
        RECT 1762.910 0.690 1766.210 4.280 ;
        RECT 1767.050 0.690 1770.350 4.280 ;
        RECT 1771.190 0.690 1774.490 4.280 ;
        RECT 1775.330 0.690 1778.630 4.280 ;
        RECT 1779.470 0.690 1782.770 4.280 ;
        RECT 1783.610 0.690 1786.910 4.280 ;
        RECT 1787.750 0.690 1791.050 4.280 ;
        RECT 1791.890 0.690 1795.190 4.280 ;
        RECT 1796.030 0.690 1799.330 4.280 ;
        RECT 1800.170 0.690 1803.470 4.280 ;
        RECT 1804.310 0.690 1807.610 4.280 ;
        RECT 1808.450 0.690 1811.750 4.280 ;
        RECT 1812.590 0.690 1815.890 4.280 ;
        RECT 1816.730 0.690 1820.030 4.280 ;
        RECT 1820.870 0.690 1824.170 4.280 ;
        RECT 1825.010 0.690 1828.310 4.280 ;
        RECT 1829.150 0.690 1832.450 4.280 ;
        RECT 1833.290 0.690 1836.590 4.280 ;
        RECT 1837.430 0.690 1840.730 4.280 ;
        RECT 1841.570 0.690 1844.870 4.280 ;
        RECT 1845.710 0.690 1849.010 4.280 ;
        RECT 1849.850 0.690 1853.150 4.280 ;
        RECT 1853.990 0.690 1857.290 4.280 ;
        RECT 1858.130 0.690 1861.430 4.280 ;
        RECT 1862.270 0.690 1865.570 4.280 ;
        RECT 1866.410 0.690 1869.710 4.280 ;
        RECT 1870.550 0.690 1873.850 4.280 ;
        RECT 1874.690 0.690 1877.990 4.280 ;
        RECT 1878.830 0.690 1882.130 4.280 ;
        RECT 1882.970 0.690 1886.270 4.280 ;
        RECT 1887.110 0.690 1890.410 4.280 ;
        RECT 1891.250 0.690 1894.550 4.280 ;
        RECT 1895.390 0.690 1898.690 4.280 ;
        RECT 1899.530 0.690 1902.830 4.280 ;
        RECT 1903.670 0.690 1906.970 4.280 ;
        RECT 1907.810 0.690 1911.110 4.280 ;
        RECT 1911.950 0.690 1915.250 4.280 ;
        RECT 1916.090 0.690 1919.390 4.280 ;
        RECT 1920.230 0.690 1923.530 4.280 ;
        RECT 1924.370 0.690 1927.670 4.280 ;
        RECT 1928.510 0.690 1931.810 4.280 ;
        RECT 1932.650 0.690 1935.950 4.280 ;
        RECT 1936.790 0.690 1940.090 4.280 ;
        RECT 1940.930 0.690 1944.230 4.280 ;
        RECT 1945.070 0.690 1948.370 4.280 ;
        RECT 1949.210 0.690 1952.510 4.280 ;
        RECT 1953.350 0.690 1956.650 4.280 ;
        RECT 1957.490 0.690 1960.790 4.280 ;
        RECT 1961.630 0.690 1964.930 4.280 ;
        RECT 1965.770 0.690 1969.070 4.280 ;
        RECT 1969.910 0.690 1973.210 4.280 ;
        RECT 1974.050 0.690 1977.350 4.280 ;
        RECT 1978.190 0.690 1981.490 4.280 ;
        RECT 1982.330 0.690 1985.630 4.280 ;
        RECT 1986.470 0.690 1989.770 4.280 ;
        RECT 1990.610 0.690 1993.910 4.280 ;
        RECT 1994.750 0.690 1998.050 4.280 ;
        RECT 1998.890 0.690 2002.190 4.280 ;
        RECT 2003.030 0.690 2006.330 4.280 ;
        RECT 2007.170 0.690 2010.470 4.280 ;
        RECT 2011.310 0.690 2014.610 4.280 ;
        RECT 2015.450 0.690 2018.750 4.280 ;
        RECT 2019.590 0.690 2022.890 4.280 ;
        RECT 2023.730 0.690 2027.030 4.280 ;
        RECT 2027.870 0.690 2031.170 4.280 ;
        RECT 2032.010 0.690 2035.310 4.280 ;
        RECT 2036.150 0.690 2039.450 4.280 ;
        RECT 2040.290 0.690 2043.590 4.280 ;
        RECT 2044.430 0.690 2047.730 4.280 ;
        RECT 2048.570 0.690 2051.870 4.280 ;
        RECT 2052.710 0.690 2056.010 4.280 ;
        RECT 2056.850 0.690 2060.150 4.280 ;
        RECT 2060.990 0.690 2064.290 4.280 ;
        RECT 2065.130 0.690 2068.430 4.280 ;
        RECT 2069.270 0.690 2072.570 4.280 ;
        RECT 2073.410 0.690 2076.710 4.280 ;
        RECT 2077.550 0.690 2080.850 4.280 ;
        RECT 2081.690 0.690 2084.990 4.280 ;
        RECT 2085.830 0.690 2089.130 4.280 ;
        RECT 2089.970 0.690 2093.270 4.280 ;
        RECT 2094.110 0.690 2097.410 4.280 ;
        RECT 2098.250 0.690 2101.550 4.280 ;
        RECT 2102.390 0.690 2105.690 4.280 ;
        RECT 2106.530 0.690 2109.830 4.280 ;
        RECT 2110.670 0.690 2113.970 4.280 ;
        RECT 2114.810 0.690 2118.110 4.280 ;
        RECT 2118.950 0.690 2195.030 4.280 ;
      LAYER met3 ;
        RECT 14.325 2.215 2195.055 2788.165 ;
      LAYER met4 ;
        RECT 15.015 10.240 20.640 2761.985 ;
        RECT 23.040 10.240 97.440 2761.985 ;
        RECT 99.840 10.240 174.240 2761.985 ;
        RECT 176.640 10.240 251.040 2761.985 ;
        RECT 253.440 10.240 327.840 2761.985 ;
        RECT 330.240 10.240 404.640 2761.985 ;
        RECT 407.040 10.240 481.440 2761.985 ;
        RECT 483.840 10.240 558.240 2761.985 ;
        RECT 560.640 10.240 635.040 2761.985 ;
        RECT 637.440 10.240 711.840 2761.985 ;
        RECT 714.240 10.240 788.640 2761.985 ;
        RECT 791.040 10.240 865.440 2761.985 ;
        RECT 867.840 10.240 942.240 2761.985 ;
        RECT 944.640 10.240 1019.040 2761.985 ;
        RECT 1021.440 10.240 1095.840 2761.985 ;
        RECT 1098.240 10.240 1172.640 2761.985 ;
        RECT 1175.040 10.240 1249.440 2761.985 ;
        RECT 1251.840 10.240 1326.240 2761.985 ;
        RECT 1328.640 10.240 1403.040 2761.985 ;
        RECT 1405.440 10.240 1479.840 2761.985 ;
        RECT 1482.240 10.240 1556.640 2761.985 ;
        RECT 1559.040 10.240 1633.440 2761.985 ;
        RECT 1635.840 10.240 1710.240 2761.985 ;
        RECT 1712.640 10.240 1787.040 2761.985 ;
        RECT 1789.440 10.240 1863.840 2761.985 ;
        RECT 1866.240 10.240 1940.640 2761.985 ;
        RECT 1943.040 10.240 2017.440 2761.985 ;
        RECT 2019.840 10.240 2094.240 2761.985 ;
        RECT 2096.640 10.240 2171.040 2761.985 ;
        RECT 2173.440 10.240 2181.025 2761.985 ;
        RECT 15.015 2.215 2181.025 10.240 ;
  END
END trainable_nn
END LIBRARY

