magic
tech sky130A
magscale 1 2
timestamp 1670254966
<< obsli1 >>
rect 1104 2159 298816 397681
<< obsm1 >>
rect 566 8 298816 397712
<< metal2 >>
rect 4434 399200 4490 400000
rect 7010 399200 7066 400000
rect 9586 399200 9642 400000
rect 12162 399200 12218 400000
rect 14738 399200 14794 400000
rect 17314 399200 17370 400000
rect 19890 399200 19946 400000
rect 22466 399200 22522 400000
rect 25042 399200 25098 400000
rect 27618 399200 27674 400000
rect 30194 399200 30250 400000
rect 32770 399200 32826 400000
rect 35346 399200 35402 400000
rect 37922 399200 37978 400000
rect 40498 399200 40554 400000
rect 43074 399200 43130 400000
rect 45650 399200 45706 400000
rect 48226 399200 48282 400000
rect 50802 399200 50858 400000
rect 53378 399200 53434 400000
rect 55954 399200 56010 400000
rect 58530 399200 58586 400000
rect 61106 399200 61162 400000
rect 63682 399200 63738 400000
rect 66258 399200 66314 400000
rect 68834 399200 68890 400000
rect 71410 399200 71466 400000
rect 73986 399200 74042 400000
rect 76562 399200 76618 400000
rect 79138 399200 79194 400000
rect 81714 399200 81770 400000
rect 84290 399200 84346 400000
rect 86866 399200 86922 400000
rect 89442 399200 89498 400000
rect 92018 399200 92074 400000
rect 94594 399200 94650 400000
rect 97170 399200 97226 400000
rect 99746 399200 99802 400000
rect 102322 399200 102378 400000
rect 104898 399200 104954 400000
rect 107474 399200 107530 400000
rect 110050 399200 110106 400000
rect 112626 399200 112682 400000
rect 115202 399200 115258 400000
rect 117778 399200 117834 400000
rect 120354 399200 120410 400000
rect 122930 399200 122986 400000
rect 125506 399200 125562 400000
rect 128082 399200 128138 400000
rect 130658 399200 130714 400000
rect 133234 399200 133290 400000
rect 135810 399200 135866 400000
rect 138386 399200 138442 400000
rect 140962 399200 141018 400000
rect 143538 399200 143594 400000
rect 146114 399200 146170 400000
rect 148690 399200 148746 400000
rect 151266 399200 151322 400000
rect 153842 399200 153898 400000
rect 156418 399200 156474 400000
rect 158994 399200 159050 400000
rect 161570 399200 161626 400000
rect 164146 399200 164202 400000
rect 166722 399200 166778 400000
rect 169298 399200 169354 400000
rect 171874 399200 171930 400000
rect 174450 399200 174506 400000
rect 177026 399200 177082 400000
rect 179602 399200 179658 400000
rect 182178 399200 182234 400000
rect 184754 399200 184810 400000
rect 187330 399200 187386 400000
rect 189906 399200 189962 400000
rect 192482 399200 192538 400000
rect 195058 399200 195114 400000
rect 197634 399200 197690 400000
rect 200210 399200 200266 400000
rect 202786 399200 202842 400000
rect 205362 399200 205418 400000
rect 207938 399200 207994 400000
rect 210514 399200 210570 400000
rect 213090 399200 213146 400000
rect 215666 399200 215722 400000
rect 218242 399200 218298 400000
rect 220818 399200 220874 400000
rect 223394 399200 223450 400000
rect 225970 399200 226026 400000
rect 228546 399200 228602 400000
rect 231122 399200 231178 400000
rect 233698 399200 233754 400000
rect 236274 399200 236330 400000
rect 238850 399200 238906 400000
rect 241426 399200 241482 400000
rect 244002 399200 244058 400000
rect 246578 399200 246634 400000
rect 249154 399200 249210 400000
rect 251730 399200 251786 400000
rect 254306 399200 254362 400000
rect 256882 399200 256938 400000
rect 259458 399200 259514 400000
rect 262034 399200 262090 400000
rect 264610 399200 264666 400000
rect 267186 399200 267242 400000
rect 269762 399200 269818 400000
rect 272338 399200 272394 400000
rect 274914 399200 274970 400000
rect 277490 399200 277546 400000
rect 280066 399200 280122 400000
rect 282642 399200 282698 400000
rect 285218 399200 285274 400000
rect 287794 399200 287850 400000
rect 290370 399200 290426 400000
rect 292946 399200 293002 400000
rect 295522 399200 295578 400000
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 60002 0 60058 800
rect 60554 0 60610 800
rect 61106 0 61162 800
rect 61658 0 61714 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65522 0 65578 800
rect 66074 0 66130 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68282 0 68338 800
rect 68834 0 68890 800
rect 69386 0 69442 800
rect 69938 0 69994 800
rect 70490 0 70546 800
rect 71042 0 71098 800
rect 71594 0 71650 800
rect 72146 0 72202 800
rect 72698 0 72754 800
rect 73250 0 73306 800
rect 73802 0 73858 800
rect 74354 0 74410 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 76010 0 76066 800
rect 76562 0 76618 800
rect 77114 0 77170 800
rect 77666 0 77722 800
rect 78218 0 78274 800
rect 78770 0 78826 800
rect 79322 0 79378 800
rect 79874 0 79930 800
rect 80426 0 80482 800
rect 80978 0 81034 800
rect 81530 0 81586 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83186 0 83242 800
rect 83738 0 83794 800
rect 84290 0 84346 800
rect 84842 0 84898 800
rect 85394 0 85450 800
rect 85946 0 86002 800
rect 86498 0 86554 800
rect 87050 0 87106 800
rect 87602 0 87658 800
rect 88154 0 88210 800
rect 88706 0 88762 800
rect 89258 0 89314 800
rect 89810 0 89866 800
rect 90362 0 90418 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93122 0 93178 800
rect 93674 0 93730 800
rect 94226 0 94282 800
rect 94778 0 94834 800
rect 95330 0 95386 800
rect 95882 0 95938 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 98090 0 98146 800
rect 98642 0 98698 800
rect 99194 0 99250 800
rect 99746 0 99802 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 101954 0 102010 800
rect 102506 0 102562 800
rect 103058 0 103114 800
rect 103610 0 103666 800
rect 104162 0 104218 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106370 0 106426 800
rect 106922 0 106978 800
rect 107474 0 107530 800
rect 108026 0 108082 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109682 0 109738 800
rect 110234 0 110290 800
rect 110786 0 110842 800
rect 111338 0 111394 800
rect 111890 0 111946 800
rect 112442 0 112498 800
rect 112994 0 113050 800
rect 113546 0 113602 800
rect 114098 0 114154 800
rect 114650 0 114706 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116306 0 116362 800
rect 116858 0 116914 800
rect 117410 0 117466 800
rect 117962 0 118018 800
rect 118514 0 118570 800
rect 119066 0 119122 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121274 0 121330 800
rect 121826 0 121882 800
rect 122378 0 122434 800
rect 122930 0 122986 800
rect 123482 0 123538 800
rect 124034 0 124090 800
rect 124586 0 124642 800
rect 125138 0 125194 800
rect 125690 0 125746 800
rect 126242 0 126298 800
rect 126794 0 126850 800
rect 127346 0 127402 800
rect 127898 0 127954 800
rect 128450 0 128506 800
rect 129002 0 129058 800
rect 129554 0 129610 800
rect 130106 0 130162 800
rect 130658 0 130714 800
rect 131210 0 131266 800
rect 131762 0 131818 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133418 0 133474 800
rect 133970 0 134026 800
rect 134522 0 134578 800
rect 135074 0 135130 800
rect 135626 0 135682 800
rect 136178 0 136234 800
rect 136730 0 136786 800
rect 137282 0 137338 800
rect 137834 0 137890 800
rect 138386 0 138442 800
rect 138938 0 138994 800
rect 139490 0 139546 800
rect 140042 0 140098 800
rect 140594 0 140650 800
rect 141146 0 141202 800
rect 141698 0 141754 800
rect 142250 0 142306 800
rect 142802 0 142858 800
rect 143354 0 143410 800
rect 143906 0 143962 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146114 0 146170 800
rect 146666 0 146722 800
rect 147218 0 147274 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148874 0 148930 800
rect 149426 0 149482 800
rect 149978 0 150034 800
rect 150530 0 150586 800
rect 151082 0 151138 800
rect 151634 0 151690 800
rect 152186 0 152242 800
rect 152738 0 152794 800
rect 153290 0 153346 800
rect 153842 0 153898 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155498 0 155554 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157154 0 157210 800
rect 157706 0 157762 800
rect 158258 0 158314 800
rect 158810 0 158866 800
rect 159362 0 159418 800
rect 159914 0 159970 800
rect 160466 0 160522 800
rect 161018 0 161074 800
rect 161570 0 161626 800
rect 162122 0 162178 800
rect 162674 0 162730 800
rect 163226 0 163282 800
rect 163778 0 163834 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 165986 0 166042 800
rect 166538 0 166594 800
rect 167090 0 167146 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168746 0 168802 800
rect 169298 0 169354 800
rect 169850 0 169906 800
rect 170402 0 170458 800
rect 170954 0 171010 800
rect 171506 0 171562 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174818 0 174874 800
rect 175370 0 175426 800
rect 175922 0 175978 800
rect 176474 0 176530 800
rect 177026 0 177082 800
rect 177578 0 177634 800
rect 178130 0 178186 800
rect 178682 0 178738 800
rect 179234 0 179290 800
rect 179786 0 179842 800
rect 180338 0 180394 800
rect 180890 0 180946 800
rect 181442 0 181498 800
rect 181994 0 182050 800
rect 182546 0 182602 800
rect 183098 0 183154 800
rect 183650 0 183706 800
rect 184202 0 184258 800
rect 184754 0 184810 800
rect 185306 0 185362 800
rect 185858 0 185914 800
rect 186410 0 186466 800
rect 186962 0 187018 800
rect 187514 0 187570 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189722 0 189778 800
rect 190274 0 190330 800
rect 190826 0 190882 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192482 0 192538 800
rect 193034 0 193090 800
rect 193586 0 193642 800
rect 194138 0 194194 800
rect 194690 0 194746 800
rect 195242 0 195298 800
rect 195794 0 195850 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197450 0 197506 800
rect 198002 0 198058 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200210 0 200266 800
rect 200762 0 200818 800
rect 201314 0 201370 800
rect 201866 0 201922 800
rect 202418 0 202474 800
rect 202970 0 203026 800
rect 203522 0 203578 800
rect 204074 0 204130 800
rect 204626 0 204682 800
rect 205178 0 205234 800
rect 205730 0 205786 800
rect 206282 0 206338 800
rect 206834 0 206890 800
rect 207386 0 207442 800
rect 207938 0 207994 800
rect 208490 0 208546 800
rect 209042 0 209098 800
rect 209594 0 209650 800
rect 210146 0 210202 800
rect 210698 0 210754 800
rect 211250 0 211306 800
rect 211802 0 211858 800
rect 212354 0 212410 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214562 0 214618 800
rect 215114 0 215170 800
rect 215666 0 215722 800
rect 216218 0 216274 800
rect 216770 0 216826 800
rect 217322 0 217378 800
rect 217874 0 217930 800
rect 218426 0 218482 800
rect 218978 0 219034 800
rect 219530 0 219586 800
rect 220082 0 220138 800
rect 220634 0 220690 800
rect 221186 0 221242 800
rect 221738 0 221794 800
rect 222290 0 222346 800
rect 222842 0 222898 800
rect 223394 0 223450 800
rect 223946 0 224002 800
rect 224498 0 224554 800
rect 225050 0 225106 800
rect 225602 0 225658 800
rect 226154 0 226210 800
rect 226706 0 226762 800
rect 227258 0 227314 800
rect 227810 0 227866 800
rect 228362 0 228418 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 230018 0 230074 800
rect 230570 0 230626 800
rect 231122 0 231178 800
rect 231674 0 231730 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233882 0 233938 800
rect 234434 0 234490 800
rect 234986 0 235042 800
rect 235538 0 235594 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237746 0 237802 800
rect 238298 0 238354 800
rect 238850 0 238906 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240506 0 240562 800
rect 241058 0 241114 800
rect 241610 0 241666 800
rect 242162 0 242218 800
rect 242714 0 242770 800
rect 243266 0 243322 800
rect 243818 0 243874 800
rect 244370 0 244426 800
rect 244922 0 244978 800
rect 245474 0 245530 800
rect 246026 0 246082 800
rect 246578 0 246634 800
rect 247130 0 247186 800
rect 247682 0 247738 800
rect 248234 0 248290 800
rect 248786 0 248842 800
rect 249338 0 249394 800
rect 249890 0 249946 800
rect 250442 0 250498 800
rect 250994 0 251050 800
rect 251546 0 251602 800
rect 252098 0 252154 800
rect 252650 0 252706 800
rect 253202 0 253258 800
rect 253754 0 253810 800
rect 254306 0 254362 800
rect 254858 0 254914 800
rect 255410 0 255466 800
rect 255962 0 256018 800
rect 256514 0 256570 800
rect 257066 0 257122 800
rect 257618 0 257674 800
rect 258170 0 258226 800
rect 258722 0 258778 800
rect 259274 0 259330 800
rect 259826 0 259882 800
rect 260378 0 260434 800
rect 260930 0 260986 800
rect 261482 0 261538 800
rect 262034 0 262090 800
rect 262586 0 262642 800
rect 263138 0 263194 800
rect 263690 0 263746 800
rect 264242 0 264298 800
rect 264794 0 264850 800
rect 265346 0 265402 800
rect 265898 0 265954 800
rect 266450 0 266506 800
rect 267002 0 267058 800
rect 267554 0 267610 800
rect 268106 0 268162 800
rect 268658 0 268714 800
rect 269210 0 269266 800
rect 269762 0 269818 800
rect 270314 0 270370 800
rect 270866 0 270922 800
rect 271418 0 271474 800
rect 271970 0 272026 800
rect 272522 0 272578 800
rect 273074 0 273130 800
rect 273626 0 273682 800
rect 274178 0 274234 800
rect 274730 0 274786 800
rect 275282 0 275338 800
rect 275834 0 275890 800
rect 276386 0 276442 800
rect 276938 0 276994 800
rect 277490 0 277546 800
rect 278042 0 278098 800
rect 278594 0 278650 800
rect 279146 0 279202 800
rect 279698 0 279754 800
rect 280250 0 280306 800
rect 280802 0 280858 800
rect 281354 0 281410 800
rect 281906 0 281962 800
rect 282458 0 282514 800
rect 283010 0 283066 800
rect 283562 0 283618 800
rect 284114 0 284170 800
rect 284666 0 284722 800
rect 285218 0 285274 800
rect 285770 0 285826 800
<< obsm2 >>
rect 570 399144 4378 399200
rect 4546 399144 6954 399200
rect 7122 399144 9530 399200
rect 9698 399144 12106 399200
rect 12274 399144 14682 399200
rect 14850 399144 17258 399200
rect 17426 399144 19834 399200
rect 20002 399144 22410 399200
rect 22578 399144 24986 399200
rect 25154 399144 27562 399200
rect 27730 399144 30138 399200
rect 30306 399144 32714 399200
rect 32882 399144 35290 399200
rect 35458 399144 37866 399200
rect 38034 399144 40442 399200
rect 40610 399144 43018 399200
rect 43186 399144 45594 399200
rect 45762 399144 48170 399200
rect 48338 399144 50746 399200
rect 50914 399144 53322 399200
rect 53490 399144 55898 399200
rect 56066 399144 58474 399200
rect 58642 399144 61050 399200
rect 61218 399144 63626 399200
rect 63794 399144 66202 399200
rect 66370 399144 68778 399200
rect 68946 399144 71354 399200
rect 71522 399144 73930 399200
rect 74098 399144 76506 399200
rect 76674 399144 79082 399200
rect 79250 399144 81658 399200
rect 81826 399144 84234 399200
rect 84402 399144 86810 399200
rect 86978 399144 89386 399200
rect 89554 399144 91962 399200
rect 92130 399144 94538 399200
rect 94706 399144 97114 399200
rect 97282 399144 99690 399200
rect 99858 399144 102266 399200
rect 102434 399144 104842 399200
rect 105010 399144 107418 399200
rect 107586 399144 109994 399200
rect 110162 399144 112570 399200
rect 112738 399144 115146 399200
rect 115314 399144 117722 399200
rect 117890 399144 120298 399200
rect 120466 399144 122874 399200
rect 123042 399144 125450 399200
rect 125618 399144 128026 399200
rect 128194 399144 130602 399200
rect 130770 399144 133178 399200
rect 133346 399144 135754 399200
rect 135922 399144 138330 399200
rect 138498 399144 140906 399200
rect 141074 399144 143482 399200
rect 143650 399144 146058 399200
rect 146226 399144 148634 399200
rect 148802 399144 151210 399200
rect 151378 399144 153786 399200
rect 153954 399144 156362 399200
rect 156530 399144 158938 399200
rect 159106 399144 161514 399200
rect 161682 399144 164090 399200
rect 164258 399144 166666 399200
rect 166834 399144 169242 399200
rect 169410 399144 171818 399200
rect 171986 399144 174394 399200
rect 174562 399144 176970 399200
rect 177138 399144 179546 399200
rect 179714 399144 182122 399200
rect 182290 399144 184698 399200
rect 184866 399144 187274 399200
rect 187442 399144 189850 399200
rect 190018 399144 192426 399200
rect 192594 399144 195002 399200
rect 195170 399144 197578 399200
rect 197746 399144 200154 399200
rect 200322 399144 202730 399200
rect 202898 399144 205306 399200
rect 205474 399144 207882 399200
rect 208050 399144 210458 399200
rect 210626 399144 213034 399200
rect 213202 399144 215610 399200
rect 215778 399144 218186 399200
rect 218354 399144 220762 399200
rect 220930 399144 223338 399200
rect 223506 399144 225914 399200
rect 226082 399144 228490 399200
rect 228658 399144 231066 399200
rect 231234 399144 233642 399200
rect 233810 399144 236218 399200
rect 236386 399144 238794 399200
rect 238962 399144 241370 399200
rect 241538 399144 243946 399200
rect 244114 399144 246522 399200
rect 246690 399144 249098 399200
rect 249266 399144 251674 399200
rect 251842 399144 254250 399200
rect 254418 399144 256826 399200
rect 256994 399144 259402 399200
rect 259570 399144 261978 399200
rect 262146 399144 264554 399200
rect 264722 399144 267130 399200
rect 267298 399144 269706 399200
rect 269874 399144 272282 399200
rect 272450 399144 274858 399200
rect 275026 399144 277434 399200
rect 277602 399144 280010 399200
rect 280178 399144 282586 399200
rect 282754 399144 285162 399200
rect 285330 399144 287738 399200
rect 287906 399144 290314 399200
rect 290482 399144 292890 399200
rect 293058 399144 295466 399200
rect 295634 399144 296362 399200
rect 570 856 296362 399144
rect 570 2 14130 856
rect 14298 2 14682 856
rect 14850 2 15234 856
rect 15402 2 15786 856
rect 15954 2 16338 856
rect 16506 2 16890 856
rect 17058 2 17442 856
rect 17610 2 17994 856
rect 18162 2 18546 856
rect 18714 2 19098 856
rect 19266 2 19650 856
rect 19818 2 20202 856
rect 20370 2 20754 856
rect 20922 2 21306 856
rect 21474 2 21858 856
rect 22026 2 22410 856
rect 22578 2 22962 856
rect 23130 2 23514 856
rect 23682 2 24066 856
rect 24234 2 24618 856
rect 24786 2 25170 856
rect 25338 2 25722 856
rect 25890 2 26274 856
rect 26442 2 26826 856
rect 26994 2 27378 856
rect 27546 2 27930 856
rect 28098 2 28482 856
rect 28650 2 29034 856
rect 29202 2 29586 856
rect 29754 2 30138 856
rect 30306 2 30690 856
rect 30858 2 31242 856
rect 31410 2 31794 856
rect 31962 2 32346 856
rect 32514 2 32898 856
rect 33066 2 33450 856
rect 33618 2 34002 856
rect 34170 2 34554 856
rect 34722 2 35106 856
rect 35274 2 35658 856
rect 35826 2 36210 856
rect 36378 2 36762 856
rect 36930 2 37314 856
rect 37482 2 37866 856
rect 38034 2 38418 856
rect 38586 2 38970 856
rect 39138 2 39522 856
rect 39690 2 40074 856
rect 40242 2 40626 856
rect 40794 2 41178 856
rect 41346 2 41730 856
rect 41898 2 42282 856
rect 42450 2 42834 856
rect 43002 2 43386 856
rect 43554 2 43938 856
rect 44106 2 44490 856
rect 44658 2 45042 856
rect 45210 2 45594 856
rect 45762 2 46146 856
rect 46314 2 46698 856
rect 46866 2 47250 856
rect 47418 2 47802 856
rect 47970 2 48354 856
rect 48522 2 48906 856
rect 49074 2 49458 856
rect 49626 2 50010 856
rect 50178 2 50562 856
rect 50730 2 51114 856
rect 51282 2 51666 856
rect 51834 2 52218 856
rect 52386 2 52770 856
rect 52938 2 53322 856
rect 53490 2 53874 856
rect 54042 2 54426 856
rect 54594 2 54978 856
rect 55146 2 55530 856
rect 55698 2 56082 856
rect 56250 2 56634 856
rect 56802 2 57186 856
rect 57354 2 57738 856
rect 57906 2 58290 856
rect 58458 2 58842 856
rect 59010 2 59394 856
rect 59562 2 59946 856
rect 60114 2 60498 856
rect 60666 2 61050 856
rect 61218 2 61602 856
rect 61770 2 62154 856
rect 62322 2 62706 856
rect 62874 2 63258 856
rect 63426 2 63810 856
rect 63978 2 64362 856
rect 64530 2 64914 856
rect 65082 2 65466 856
rect 65634 2 66018 856
rect 66186 2 66570 856
rect 66738 2 67122 856
rect 67290 2 67674 856
rect 67842 2 68226 856
rect 68394 2 68778 856
rect 68946 2 69330 856
rect 69498 2 69882 856
rect 70050 2 70434 856
rect 70602 2 70986 856
rect 71154 2 71538 856
rect 71706 2 72090 856
rect 72258 2 72642 856
rect 72810 2 73194 856
rect 73362 2 73746 856
rect 73914 2 74298 856
rect 74466 2 74850 856
rect 75018 2 75402 856
rect 75570 2 75954 856
rect 76122 2 76506 856
rect 76674 2 77058 856
rect 77226 2 77610 856
rect 77778 2 78162 856
rect 78330 2 78714 856
rect 78882 2 79266 856
rect 79434 2 79818 856
rect 79986 2 80370 856
rect 80538 2 80922 856
rect 81090 2 81474 856
rect 81642 2 82026 856
rect 82194 2 82578 856
rect 82746 2 83130 856
rect 83298 2 83682 856
rect 83850 2 84234 856
rect 84402 2 84786 856
rect 84954 2 85338 856
rect 85506 2 85890 856
rect 86058 2 86442 856
rect 86610 2 86994 856
rect 87162 2 87546 856
rect 87714 2 88098 856
rect 88266 2 88650 856
rect 88818 2 89202 856
rect 89370 2 89754 856
rect 89922 2 90306 856
rect 90474 2 90858 856
rect 91026 2 91410 856
rect 91578 2 91962 856
rect 92130 2 92514 856
rect 92682 2 93066 856
rect 93234 2 93618 856
rect 93786 2 94170 856
rect 94338 2 94722 856
rect 94890 2 95274 856
rect 95442 2 95826 856
rect 95994 2 96378 856
rect 96546 2 96930 856
rect 97098 2 97482 856
rect 97650 2 98034 856
rect 98202 2 98586 856
rect 98754 2 99138 856
rect 99306 2 99690 856
rect 99858 2 100242 856
rect 100410 2 100794 856
rect 100962 2 101346 856
rect 101514 2 101898 856
rect 102066 2 102450 856
rect 102618 2 103002 856
rect 103170 2 103554 856
rect 103722 2 104106 856
rect 104274 2 104658 856
rect 104826 2 105210 856
rect 105378 2 105762 856
rect 105930 2 106314 856
rect 106482 2 106866 856
rect 107034 2 107418 856
rect 107586 2 107970 856
rect 108138 2 108522 856
rect 108690 2 109074 856
rect 109242 2 109626 856
rect 109794 2 110178 856
rect 110346 2 110730 856
rect 110898 2 111282 856
rect 111450 2 111834 856
rect 112002 2 112386 856
rect 112554 2 112938 856
rect 113106 2 113490 856
rect 113658 2 114042 856
rect 114210 2 114594 856
rect 114762 2 115146 856
rect 115314 2 115698 856
rect 115866 2 116250 856
rect 116418 2 116802 856
rect 116970 2 117354 856
rect 117522 2 117906 856
rect 118074 2 118458 856
rect 118626 2 119010 856
rect 119178 2 119562 856
rect 119730 2 120114 856
rect 120282 2 120666 856
rect 120834 2 121218 856
rect 121386 2 121770 856
rect 121938 2 122322 856
rect 122490 2 122874 856
rect 123042 2 123426 856
rect 123594 2 123978 856
rect 124146 2 124530 856
rect 124698 2 125082 856
rect 125250 2 125634 856
rect 125802 2 126186 856
rect 126354 2 126738 856
rect 126906 2 127290 856
rect 127458 2 127842 856
rect 128010 2 128394 856
rect 128562 2 128946 856
rect 129114 2 129498 856
rect 129666 2 130050 856
rect 130218 2 130602 856
rect 130770 2 131154 856
rect 131322 2 131706 856
rect 131874 2 132258 856
rect 132426 2 132810 856
rect 132978 2 133362 856
rect 133530 2 133914 856
rect 134082 2 134466 856
rect 134634 2 135018 856
rect 135186 2 135570 856
rect 135738 2 136122 856
rect 136290 2 136674 856
rect 136842 2 137226 856
rect 137394 2 137778 856
rect 137946 2 138330 856
rect 138498 2 138882 856
rect 139050 2 139434 856
rect 139602 2 139986 856
rect 140154 2 140538 856
rect 140706 2 141090 856
rect 141258 2 141642 856
rect 141810 2 142194 856
rect 142362 2 142746 856
rect 142914 2 143298 856
rect 143466 2 143850 856
rect 144018 2 144402 856
rect 144570 2 144954 856
rect 145122 2 145506 856
rect 145674 2 146058 856
rect 146226 2 146610 856
rect 146778 2 147162 856
rect 147330 2 147714 856
rect 147882 2 148266 856
rect 148434 2 148818 856
rect 148986 2 149370 856
rect 149538 2 149922 856
rect 150090 2 150474 856
rect 150642 2 151026 856
rect 151194 2 151578 856
rect 151746 2 152130 856
rect 152298 2 152682 856
rect 152850 2 153234 856
rect 153402 2 153786 856
rect 153954 2 154338 856
rect 154506 2 154890 856
rect 155058 2 155442 856
rect 155610 2 155994 856
rect 156162 2 156546 856
rect 156714 2 157098 856
rect 157266 2 157650 856
rect 157818 2 158202 856
rect 158370 2 158754 856
rect 158922 2 159306 856
rect 159474 2 159858 856
rect 160026 2 160410 856
rect 160578 2 160962 856
rect 161130 2 161514 856
rect 161682 2 162066 856
rect 162234 2 162618 856
rect 162786 2 163170 856
rect 163338 2 163722 856
rect 163890 2 164274 856
rect 164442 2 164826 856
rect 164994 2 165378 856
rect 165546 2 165930 856
rect 166098 2 166482 856
rect 166650 2 167034 856
rect 167202 2 167586 856
rect 167754 2 168138 856
rect 168306 2 168690 856
rect 168858 2 169242 856
rect 169410 2 169794 856
rect 169962 2 170346 856
rect 170514 2 170898 856
rect 171066 2 171450 856
rect 171618 2 172002 856
rect 172170 2 172554 856
rect 172722 2 173106 856
rect 173274 2 173658 856
rect 173826 2 174210 856
rect 174378 2 174762 856
rect 174930 2 175314 856
rect 175482 2 175866 856
rect 176034 2 176418 856
rect 176586 2 176970 856
rect 177138 2 177522 856
rect 177690 2 178074 856
rect 178242 2 178626 856
rect 178794 2 179178 856
rect 179346 2 179730 856
rect 179898 2 180282 856
rect 180450 2 180834 856
rect 181002 2 181386 856
rect 181554 2 181938 856
rect 182106 2 182490 856
rect 182658 2 183042 856
rect 183210 2 183594 856
rect 183762 2 184146 856
rect 184314 2 184698 856
rect 184866 2 185250 856
rect 185418 2 185802 856
rect 185970 2 186354 856
rect 186522 2 186906 856
rect 187074 2 187458 856
rect 187626 2 188010 856
rect 188178 2 188562 856
rect 188730 2 189114 856
rect 189282 2 189666 856
rect 189834 2 190218 856
rect 190386 2 190770 856
rect 190938 2 191322 856
rect 191490 2 191874 856
rect 192042 2 192426 856
rect 192594 2 192978 856
rect 193146 2 193530 856
rect 193698 2 194082 856
rect 194250 2 194634 856
rect 194802 2 195186 856
rect 195354 2 195738 856
rect 195906 2 196290 856
rect 196458 2 196842 856
rect 197010 2 197394 856
rect 197562 2 197946 856
rect 198114 2 198498 856
rect 198666 2 199050 856
rect 199218 2 199602 856
rect 199770 2 200154 856
rect 200322 2 200706 856
rect 200874 2 201258 856
rect 201426 2 201810 856
rect 201978 2 202362 856
rect 202530 2 202914 856
rect 203082 2 203466 856
rect 203634 2 204018 856
rect 204186 2 204570 856
rect 204738 2 205122 856
rect 205290 2 205674 856
rect 205842 2 206226 856
rect 206394 2 206778 856
rect 206946 2 207330 856
rect 207498 2 207882 856
rect 208050 2 208434 856
rect 208602 2 208986 856
rect 209154 2 209538 856
rect 209706 2 210090 856
rect 210258 2 210642 856
rect 210810 2 211194 856
rect 211362 2 211746 856
rect 211914 2 212298 856
rect 212466 2 212850 856
rect 213018 2 213402 856
rect 213570 2 213954 856
rect 214122 2 214506 856
rect 214674 2 215058 856
rect 215226 2 215610 856
rect 215778 2 216162 856
rect 216330 2 216714 856
rect 216882 2 217266 856
rect 217434 2 217818 856
rect 217986 2 218370 856
rect 218538 2 218922 856
rect 219090 2 219474 856
rect 219642 2 220026 856
rect 220194 2 220578 856
rect 220746 2 221130 856
rect 221298 2 221682 856
rect 221850 2 222234 856
rect 222402 2 222786 856
rect 222954 2 223338 856
rect 223506 2 223890 856
rect 224058 2 224442 856
rect 224610 2 224994 856
rect 225162 2 225546 856
rect 225714 2 226098 856
rect 226266 2 226650 856
rect 226818 2 227202 856
rect 227370 2 227754 856
rect 227922 2 228306 856
rect 228474 2 228858 856
rect 229026 2 229410 856
rect 229578 2 229962 856
rect 230130 2 230514 856
rect 230682 2 231066 856
rect 231234 2 231618 856
rect 231786 2 232170 856
rect 232338 2 232722 856
rect 232890 2 233274 856
rect 233442 2 233826 856
rect 233994 2 234378 856
rect 234546 2 234930 856
rect 235098 2 235482 856
rect 235650 2 236034 856
rect 236202 2 236586 856
rect 236754 2 237138 856
rect 237306 2 237690 856
rect 237858 2 238242 856
rect 238410 2 238794 856
rect 238962 2 239346 856
rect 239514 2 239898 856
rect 240066 2 240450 856
rect 240618 2 241002 856
rect 241170 2 241554 856
rect 241722 2 242106 856
rect 242274 2 242658 856
rect 242826 2 243210 856
rect 243378 2 243762 856
rect 243930 2 244314 856
rect 244482 2 244866 856
rect 245034 2 245418 856
rect 245586 2 245970 856
rect 246138 2 246522 856
rect 246690 2 247074 856
rect 247242 2 247626 856
rect 247794 2 248178 856
rect 248346 2 248730 856
rect 248898 2 249282 856
rect 249450 2 249834 856
rect 250002 2 250386 856
rect 250554 2 250938 856
rect 251106 2 251490 856
rect 251658 2 252042 856
rect 252210 2 252594 856
rect 252762 2 253146 856
rect 253314 2 253698 856
rect 253866 2 254250 856
rect 254418 2 254802 856
rect 254970 2 255354 856
rect 255522 2 255906 856
rect 256074 2 256458 856
rect 256626 2 257010 856
rect 257178 2 257562 856
rect 257730 2 258114 856
rect 258282 2 258666 856
rect 258834 2 259218 856
rect 259386 2 259770 856
rect 259938 2 260322 856
rect 260490 2 260874 856
rect 261042 2 261426 856
rect 261594 2 261978 856
rect 262146 2 262530 856
rect 262698 2 263082 856
rect 263250 2 263634 856
rect 263802 2 264186 856
rect 264354 2 264738 856
rect 264906 2 265290 856
rect 265458 2 265842 856
rect 266010 2 266394 856
rect 266562 2 266946 856
rect 267114 2 267498 856
rect 267666 2 268050 856
rect 268218 2 268602 856
rect 268770 2 269154 856
rect 269322 2 269706 856
rect 269874 2 270258 856
rect 270426 2 270810 856
rect 270978 2 271362 856
rect 271530 2 271914 856
rect 272082 2 272466 856
rect 272634 2 273018 856
rect 273186 2 273570 856
rect 273738 2 274122 856
rect 274290 2 274674 856
rect 274842 2 275226 856
rect 275394 2 275778 856
rect 275946 2 276330 856
rect 276498 2 276882 856
rect 277050 2 277434 856
rect 277602 2 277986 856
rect 278154 2 278538 856
rect 278706 2 279090 856
rect 279258 2 279642 856
rect 279810 2 280194 856
rect 280362 2 280746 856
rect 280914 2 281298 856
rect 281466 2 281850 856
rect 282018 2 282402 856
rect 282570 2 282954 856
rect 283122 2 283506 856
rect 283674 2 284058 856
rect 284226 2 284610 856
rect 284778 2 285162 856
rect 285330 2 285714 856
rect 285882 2 296362 856
<< obsm3 >>
rect 565 443 296366 397697
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
rect 203888 2128 204208 397712
rect 219248 2128 219568 397712
rect 234608 2128 234928 397712
rect 249968 2128 250288 397712
rect 265328 2128 265648 397712
rect 280688 2128 281008 397712
rect 296048 2128 296368 397712
<< obsm4 >>
rect 979 2048 4128 390829
rect 4608 2048 19488 390829
rect 19968 2048 34848 390829
rect 35328 2048 50208 390829
rect 50688 2048 65568 390829
rect 66048 2048 80928 390829
rect 81408 2048 96288 390829
rect 96768 2048 111648 390829
rect 112128 2048 127008 390829
rect 127488 2048 142368 390829
rect 142848 2048 157728 390829
rect 158208 2048 173088 390829
rect 173568 2048 188448 390829
rect 188928 2048 203808 390829
rect 204288 2048 219168 390829
rect 219648 2048 234528 390829
rect 235008 2048 249888 390829
rect 250368 2048 265248 390829
rect 265728 2048 280608 390829
rect 281088 2048 290109 390829
rect 979 443 290109 2048
<< labels >>
rlabel metal2 s 4434 399200 4490 400000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 81714 399200 81770 400000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 89442 399200 89498 400000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 97170 399200 97226 400000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 104898 399200 104954 400000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 112626 399200 112682 400000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 120354 399200 120410 400000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 128082 399200 128138 400000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 135810 399200 135866 400000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 143538 399200 143594 400000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 151266 399200 151322 400000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12162 399200 12218 400000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 158994 399200 159050 400000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 166722 399200 166778 400000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 174450 399200 174506 400000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 182178 399200 182234 400000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 189906 399200 189962 400000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 197634 399200 197690 400000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 205362 399200 205418 400000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 213090 399200 213146 400000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 220818 399200 220874 400000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 228546 399200 228602 400000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 19890 399200 19946 400000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 236274 399200 236330 400000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 244002 399200 244058 400000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 251730 399200 251786 400000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 259458 399200 259514 400000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 267186 399200 267242 400000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 274914 399200 274970 400000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 282642 399200 282698 400000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 290370 399200 290426 400000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 27618 399200 27674 400000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 35346 399200 35402 400000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 43074 399200 43130 400000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 50802 399200 50858 400000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 58530 399200 58586 400000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 66258 399200 66314 400000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 73986 399200 74042 400000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 7010 399200 7066 400000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 84290 399200 84346 400000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 92018 399200 92074 400000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 99746 399200 99802 400000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 107474 399200 107530 400000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 115202 399200 115258 400000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 122930 399200 122986 400000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 130658 399200 130714 400000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 138386 399200 138442 400000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 146114 399200 146170 400000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 153842 399200 153898 400000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 14738 399200 14794 400000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 161570 399200 161626 400000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 169298 399200 169354 400000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 177026 399200 177082 400000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 184754 399200 184810 400000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 192482 399200 192538 400000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 200210 399200 200266 400000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 207938 399200 207994 400000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 215666 399200 215722 400000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 223394 399200 223450 400000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 231122 399200 231178 400000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 22466 399200 22522 400000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 238850 399200 238906 400000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 246578 399200 246634 400000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 254306 399200 254362 400000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 262034 399200 262090 400000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 269762 399200 269818 400000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 277490 399200 277546 400000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 285218 399200 285274 400000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 292946 399200 293002 400000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 30194 399200 30250 400000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 37922 399200 37978 400000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 45650 399200 45706 400000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 53378 399200 53434 400000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 61106 399200 61162 400000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 68834 399200 68890 400000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 76562 399200 76618 400000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9586 399200 9642 400000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 86866 399200 86922 400000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 94594 399200 94650 400000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 102322 399200 102378 400000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 110050 399200 110106 400000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 117778 399200 117834 400000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 125506 399200 125562 400000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 133234 399200 133290 400000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 140962 399200 141018 400000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 148690 399200 148746 400000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 156418 399200 156474 400000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 17314 399200 17370 400000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 164146 399200 164202 400000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 171874 399200 171930 400000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 179602 399200 179658 400000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 187330 399200 187386 400000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 195058 399200 195114 400000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 202786 399200 202842 400000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 210514 399200 210570 400000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 218242 399200 218298 400000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 225970 399200 226026 400000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 233698 399200 233754 400000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 25042 399200 25098 400000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 241426 399200 241482 400000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 249154 399200 249210 400000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 256882 399200 256938 400000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 264610 399200 264666 400000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 272338 399200 272394 400000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 280066 399200 280122 400000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 287794 399200 287850 400000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 295522 399200 295578 400000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 32770 399200 32826 400000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 40498 399200 40554 400000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 48226 399200 48282 400000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 55954 399200 56010 400000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 63682 399200 63738 400000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 71410 399200 71466 400000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 79138 399200 79194 400000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 284666 0 284722 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 285218 0 285274 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 285770 0 285826 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 238298 0 238354 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 241610 0 241666 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 251546 0 251602 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 253202 0 253258 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 256514 0 256570 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 269762 0 269818 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 271418 0 271474 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 276386 0 276442 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 278042 0 278098 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 279698 0 279754 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 206834 0 206890 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 216770 0 216826 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 231674 0 231730 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 238850 0 238906 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 243818 0 243874 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 245474 0 245530 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 247130 0 247186 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 248786 0 248842 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 250442 0 250498 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 252098 0 252154 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 255410 0 255466 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 258722 0 258778 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 260378 0 260434 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 263690 0 263746 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 265346 0 265402 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 267002 0 267058 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 268658 0 268714 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 270314 0 270370 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 271970 0 272026 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 273626 0 273682 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 275282 0 275338 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 276938 0 276994 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 278594 0 278650 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 280250 0 280306 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 170954 0 171010 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 174266 0 174322 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 179234 0 179290 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 182546 0 182602 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 189170 0 189226 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 200762 0 200818 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 205730 0 205786 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 207386 0 207442 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 209042 0 209098 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 210698 0 210754 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 212354 0 212410 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 214010 0 214066 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 220634 0 220690 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 222290 0 222346 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 225602 0 225658 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 227258 0 227314 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 230570 0 230626 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 235538 0 235594 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 237194 0 237250 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 241058 0 241114 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 247682 0 247738 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 249338 0 249394 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 250994 0 251050 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 260930 0 260986 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 262586 0 262642 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 274178 0 274234 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 277490 0 277546 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 279146 0 279202 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 282458 0 282514 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 201314 0 201370 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 202970 0 203026 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 207938 0 207994 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 219530 0 219586 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 227810 0 227866 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 397712 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 397712 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 14186 0 14242 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 400000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 370794980
string GDS_FILE /home/htamas/progs/trainable-nn-resub4/openlane/trainable_nn/runs/22_12_05_11_34/results/signoff/trainable_nn.magic.gds
string GDS_START 1866478
<< end >>

