magic
tech sky130B
magscale 1 2
timestamp 1657064826
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 756 178848 117552
<< metal2 >>
rect 1582 119200 1638 120000
rect 3146 119200 3202 120000
rect 4710 119200 4766 120000
rect 6274 119200 6330 120000
rect 7838 119200 7894 120000
rect 9402 119200 9458 120000
rect 10966 119200 11022 120000
rect 12530 119200 12586 120000
rect 14094 119200 14150 120000
rect 15658 119200 15714 120000
rect 17222 119200 17278 120000
rect 18786 119200 18842 120000
rect 20350 119200 20406 120000
rect 21914 119200 21970 120000
rect 23478 119200 23534 120000
rect 25042 119200 25098 120000
rect 26606 119200 26662 120000
rect 28170 119200 28226 120000
rect 29734 119200 29790 120000
rect 31298 119200 31354 120000
rect 32862 119200 32918 120000
rect 34426 119200 34482 120000
rect 35990 119200 36046 120000
rect 37554 119200 37610 120000
rect 39118 119200 39174 120000
rect 40682 119200 40738 120000
rect 42246 119200 42302 120000
rect 43810 119200 43866 120000
rect 45374 119200 45430 120000
rect 46938 119200 46994 120000
rect 48502 119200 48558 120000
rect 50066 119200 50122 120000
rect 51630 119200 51686 120000
rect 53194 119200 53250 120000
rect 54758 119200 54814 120000
rect 56322 119200 56378 120000
rect 57886 119200 57942 120000
rect 59450 119200 59506 120000
rect 61014 119200 61070 120000
rect 62578 119200 62634 120000
rect 64142 119200 64198 120000
rect 65706 119200 65762 120000
rect 67270 119200 67326 120000
rect 68834 119200 68890 120000
rect 70398 119200 70454 120000
rect 71962 119200 72018 120000
rect 73526 119200 73582 120000
rect 75090 119200 75146 120000
rect 76654 119200 76710 120000
rect 78218 119200 78274 120000
rect 79782 119200 79838 120000
rect 81346 119200 81402 120000
rect 82910 119200 82966 120000
rect 84474 119200 84530 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95422 119200 95478 120000
rect 96986 119200 97042 120000
rect 98550 119200 98606 120000
rect 100114 119200 100170 120000
rect 101678 119200 101734 120000
rect 103242 119200 103298 120000
rect 104806 119200 104862 120000
rect 106370 119200 106426 120000
rect 107934 119200 107990 120000
rect 109498 119200 109554 120000
rect 111062 119200 111118 120000
rect 112626 119200 112682 120000
rect 114190 119200 114246 120000
rect 115754 119200 115810 120000
rect 117318 119200 117374 120000
rect 118882 119200 118938 120000
rect 120446 119200 120502 120000
rect 122010 119200 122066 120000
rect 123574 119200 123630 120000
rect 125138 119200 125194 120000
rect 126702 119200 126758 120000
rect 128266 119200 128322 120000
rect 129830 119200 129886 120000
rect 131394 119200 131450 120000
rect 132958 119200 133014 120000
rect 134522 119200 134578 120000
rect 136086 119200 136142 120000
rect 137650 119200 137706 120000
rect 139214 119200 139270 120000
rect 140778 119200 140834 120000
rect 142342 119200 142398 120000
rect 143906 119200 143962 120000
rect 145470 119200 145526 120000
rect 147034 119200 147090 120000
rect 148598 119200 148654 120000
rect 150162 119200 150218 120000
rect 151726 119200 151782 120000
rect 153290 119200 153346 120000
rect 154854 119200 154910 120000
rect 156418 119200 156474 120000
rect 157982 119200 158038 120000
rect 159546 119200 159602 120000
rect 161110 119200 161166 120000
rect 162674 119200 162730 120000
rect 164238 119200 164294 120000
rect 165802 119200 165858 120000
rect 167366 119200 167422 120000
rect 168930 119200 168986 120000
rect 170494 119200 170550 120000
rect 172058 119200 172114 120000
rect 173622 119200 173678 120000
rect 175186 119200 175242 120000
rect 176750 119200 176806 120000
rect 178314 119200 178370 120000
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 38934 0 38990 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 46938 0 46994 800
rect 47214 0 47270 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54114 0 54170 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64878 0 64934 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67086 0 67142 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68742 0 68798 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72606 0 72662 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 75090 0 75146 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84198 0 84254 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94686 0 94742 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98550 0 98606 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102138 0 102194 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 106002 0 106058 800
rect 106278 0 106334 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109038 0 109094 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110142 0 110198 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114558 0 114614 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115938 0 115994 800
rect 116214 0 116270 800
rect 116490 0 116546 800
rect 116766 0 116822 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120078 0 120134 800
rect 120354 0 120410 800
rect 120630 0 120686 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123114 0 123170 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 123942 0 123998 800
rect 124218 0 124274 800
rect 124494 0 124550 800
rect 124770 0 124826 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125598 0 125654 800
rect 125874 0 125930 800
rect 126150 0 126206 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128634 0 128690 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130290 0 130346 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131118 0 131174 800
rect 131394 0 131450 800
rect 131670 0 131726 800
rect 131946 0 132002 800
rect 132222 0 132278 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134154 0 134210 800
rect 134430 0 134486 800
rect 134706 0 134762 800
rect 134982 0 135038 800
rect 135258 0 135314 800
rect 135534 0 135590 800
rect 135810 0 135866 800
rect 136086 0 136142 800
rect 136362 0 136418 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137190 0 137246 800
rect 137466 0 137522 800
rect 137742 0 137798 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139122 0 139178 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140502 0 140558 800
rect 140778 0 140834 800
rect 141054 0 141110 800
rect 141330 0 141386 800
rect 141606 0 141662 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142434 0 142490 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144090 0 144146 800
rect 144366 0 144422 800
rect 144642 0 144698 800
rect 144918 0 144974 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146022 0 146078 800
rect 146298 0 146354 800
rect 146574 0 146630 800
rect 146850 0 146906 800
rect 147126 0 147182 800
rect 147402 0 147458 800
rect 147678 0 147734 800
rect 147954 0 148010 800
rect 148230 0 148286 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149610 0 149666 800
rect 149886 0 149942 800
rect 150162 0 150218 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 150990 0 151046 800
rect 151266 0 151322 800
rect 151542 0 151598 800
rect 151818 0 151874 800
rect 152094 0 152150 800
rect 152370 0 152426 800
rect 152646 0 152702 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153474 0 153530 800
rect 153750 0 153806 800
rect 154026 0 154082 800
rect 154302 0 154358 800
rect 154578 0 154634 800
rect 154854 0 154910 800
rect 155130 0 155186 800
rect 155406 0 155462 800
rect 155682 0 155738 800
rect 155958 0 156014 800
rect 156234 0 156290 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157062 0 157118 800
rect 157338 0 157394 800
rect 157614 0 157670 800
rect 157890 0 157946 800
<< obsm2 >>
rect 3258 119144 4654 119354
rect 4822 119144 6218 119354
rect 6386 119144 7782 119354
rect 7950 119144 9346 119354
rect 9514 119144 10910 119354
rect 11078 119144 12474 119354
rect 12642 119144 14038 119354
rect 14206 119144 15602 119354
rect 15770 119144 17166 119354
rect 17334 119144 18730 119354
rect 18898 119144 20294 119354
rect 20462 119144 21858 119354
rect 22026 119144 23422 119354
rect 23590 119144 24986 119354
rect 25154 119144 26550 119354
rect 26718 119144 28114 119354
rect 28282 119144 29678 119354
rect 29846 119144 31242 119354
rect 31410 119144 32806 119354
rect 32974 119144 34370 119354
rect 34538 119144 35934 119354
rect 36102 119144 37498 119354
rect 37666 119144 39062 119354
rect 39230 119144 40626 119354
rect 40794 119144 42190 119354
rect 42358 119144 43754 119354
rect 43922 119144 45318 119354
rect 45486 119144 46882 119354
rect 47050 119144 48446 119354
rect 48614 119144 50010 119354
rect 50178 119144 51574 119354
rect 51742 119144 53138 119354
rect 53306 119144 54702 119354
rect 54870 119144 56266 119354
rect 56434 119144 57830 119354
rect 57998 119144 59394 119354
rect 59562 119144 60958 119354
rect 61126 119144 62522 119354
rect 62690 119144 64086 119354
rect 64254 119144 65650 119354
rect 65818 119144 67214 119354
rect 67382 119144 68778 119354
rect 68946 119144 70342 119354
rect 70510 119144 71906 119354
rect 72074 119144 73470 119354
rect 73638 119144 75034 119354
rect 75202 119144 76598 119354
rect 76766 119144 78162 119354
rect 78330 119144 79726 119354
rect 79894 119144 81290 119354
rect 81458 119144 82854 119354
rect 83022 119144 84418 119354
rect 84586 119144 85982 119354
rect 86150 119144 87546 119354
rect 87714 119144 89110 119354
rect 89278 119144 90674 119354
rect 90842 119144 92238 119354
rect 92406 119144 93802 119354
rect 93970 119144 95366 119354
rect 95534 119144 96930 119354
rect 97098 119144 98494 119354
rect 98662 119144 100058 119354
rect 100226 119144 101622 119354
rect 101790 119144 103186 119354
rect 103354 119144 104750 119354
rect 104918 119144 106314 119354
rect 106482 119144 107878 119354
rect 108046 119144 109442 119354
rect 109610 119144 111006 119354
rect 111174 119144 112570 119354
rect 112738 119144 114134 119354
rect 114302 119144 115698 119354
rect 115866 119144 117262 119354
rect 117430 119144 118826 119354
rect 118994 119144 120390 119354
rect 120558 119144 121954 119354
rect 122122 119144 123518 119354
rect 123686 119144 125082 119354
rect 125250 119144 126646 119354
rect 126814 119144 128210 119354
rect 128378 119144 129774 119354
rect 129942 119144 131338 119354
rect 131506 119144 132902 119354
rect 133070 119144 134466 119354
rect 134634 119144 136030 119354
rect 136198 119144 137594 119354
rect 137762 119144 139158 119354
rect 139326 119144 140722 119354
rect 140890 119144 142286 119354
rect 142454 119144 143850 119354
rect 144018 119144 145414 119354
rect 145582 119144 146978 119354
rect 147146 119144 148542 119354
rect 148710 119144 150106 119354
rect 150274 119144 151670 119354
rect 151838 119144 153234 119354
rect 153402 119144 154798 119354
rect 154966 119144 156362 119354
rect 156530 119144 157926 119354
rect 158094 119144 159490 119354
rect 159658 119144 161054 119354
rect 161222 119144 162618 119354
rect 162786 119144 164182 119354
rect 164350 119144 165746 119354
rect 165914 119144 167310 119354
rect 167478 119144 168874 119354
rect 169042 119144 170438 119354
rect 170606 119144 172002 119354
rect 172170 119144 173566 119354
rect 173734 119144 175130 119354
rect 175298 119144 176694 119354
rect 176862 119144 178258 119354
rect 3148 856 178314 119144
rect 3148 734 22042 856
rect 22210 734 22318 856
rect 22486 734 22594 856
rect 22762 734 22870 856
rect 23038 734 23146 856
rect 23314 734 23422 856
rect 23590 734 23698 856
rect 23866 734 23974 856
rect 24142 734 24250 856
rect 24418 734 24526 856
rect 24694 734 24802 856
rect 24970 734 25078 856
rect 25246 734 25354 856
rect 25522 734 25630 856
rect 25798 734 25906 856
rect 26074 734 26182 856
rect 26350 734 26458 856
rect 26626 734 26734 856
rect 26902 734 27010 856
rect 27178 734 27286 856
rect 27454 734 27562 856
rect 27730 734 27838 856
rect 28006 734 28114 856
rect 28282 734 28390 856
rect 28558 734 28666 856
rect 28834 734 28942 856
rect 29110 734 29218 856
rect 29386 734 29494 856
rect 29662 734 29770 856
rect 29938 734 30046 856
rect 30214 734 30322 856
rect 30490 734 30598 856
rect 30766 734 30874 856
rect 31042 734 31150 856
rect 31318 734 31426 856
rect 31594 734 31702 856
rect 31870 734 31978 856
rect 32146 734 32254 856
rect 32422 734 32530 856
rect 32698 734 32806 856
rect 32974 734 33082 856
rect 33250 734 33358 856
rect 33526 734 33634 856
rect 33802 734 33910 856
rect 34078 734 34186 856
rect 34354 734 34462 856
rect 34630 734 34738 856
rect 34906 734 35014 856
rect 35182 734 35290 856
rect 35458 734 35566 856
rect 35734 734 35842 856
rect 36010 734 36118 856
rect 36286 734 36394 856
rect 36562 734 36670 856
rect 36838 734 36946 856
rect 37114 734 37222 856
rect 37390 734 37498 856
rect 37666 734 37774 856
rect 37942 734 38050 856
rect 38218 734 38326 856
rect 38494 734 38602 856
rect 38770 734 38878 856
rect 39046 734 39154 856
rect 39322 734 39430 856
rect 39598 734 39706 856
rect 39874 734 39982 856
rect 40150 734 40258 856
rect 40426 734 40534 856
rect 40702 734 40810 856
rect 40978 734 41086 856
rect 41254 734 41362 856
rect 41530 734 41638 856
rect 41806 734 41914 856
rect 42082 734 42190 856
rect 42358 734 42466 856
rect 42634 734 42742 856
rect 42910 734 43018 856
rect 43186 734 43294 856
rect 43462 734 43570 856
rect 43738 734 43846 856
rect 44014 734 44122 856
rect 44290 734 44398 856
rect 44566 734 44674 856
rect 44842 734 44950 856
rect 45118 734 45226 856
rect 45394 734 45502 856
rect 45670 734 45778 856
rect 45946 734 46054 856
rect 46222 734 46330 856
rect 46498 734 46606 856
rect 46774 734 46882 856
rect 47050 734 47158 856
rect 47326 734 47434 856
rect 47602 734 47710 856
rect 47878 734 47986 856
rect 48154 734 48262 856
rect 48430 734 48538 856
rect 48706 734 48814 856
rect 48982 734 49090 856
rect 49258 734 49366 856
rect 49534 734 49642 856
rect 49810 734 49918 856
rect 50086 734 50194 856
rect 50362 734 50470 856
rect 50638 734 50746 856
rect 50914 734 51022 856
rect 51190 734 51298 856
rect 51466 734 51574 856
rect 51742 734 51850 856
rect 52018 734 52126 856
rect 52294 734 52402 856
rect 52570 734 52678 856
rect 52846 734 52954 856
rect 53122 734 53230 856
rect 53398 734 53506 856
rect 53674 734 53782 856
rect 53950 734 54058 856
rect 54226 734 54334 856
rect 54502 734 54610 856
rect 54778 734 54886 856
rect 55054 734 55162 856
rect 55330 734 55438 856
rect 55606 734 55714 856
rect 55882 734 55990 856
rect 56158 734 56266 856
rect 56434 734 56542 856
rect 56710 734 56818 856
rect 56986 734 57094 856
rect 57262 734 57370 856
rect 57538 734 57646 856
rect 57814 734 57922 856
rect 58090 734 58198 856
rect 58366 734 58474 856
rect 58642 734 58750 856
rect 58918 734 59026 856
rect 59194 734 59302 856
rect 59470 734 59578 856
rect 59746 734 59854 856
rect 60022 734 60130 856
rect 60298 734 60406 856
rect 60574 734 60682 856
rect 60850 734 60958 856
rect 61126 734 61234 856
rect 61402 734 61510 856
rect 61678 734 61786 856
rect 61954 734 62062 856
rect 62230 734 62338 856
rect 62506 734 62614 856
rect 62782 734 62890 856
rect 63058 734 63166 856
rect 63334 734 63442 856
rect 63610 734 63718 856
rect 63886 734 63994 856
rect 64162 734 64270 856
rect 64438 734 64546 856
rect 64714 734 64822 856
rect 64990 734 65098 856
rect 65266 734 65374 856
rect 65542 734 65650 856
rect 65818 734 65926 856
rect 66094 734 66202 856
rect 66370 734 66478 856
rect 66646 734 66754 856
rect 66922 734 67030 856
rect 67198 734 67306 856
rect 67474 734 67582 856
rect 67750 734 67858 856
rect 68026 734 68134 856
rect 68302 734 68410 856
rect 68578 734 68686 856
rect 68854 734 68962 856
rect 69130 734 69238 856
rect 69406 734 69514 856
rect 69682 734 69790 856
rect 69958 734 70066 856
rect 70234 734 70342 856
rect 70510 734 70618 856
rect 70786 734 70894 856
rect 71062 734 71170 856
rect 71338 734 71446 856
rect 71614 734 71722 856
rect 71890 734 71998 856
rect 72166 734 72274 856
rect 72442 734 72550 856
rect 72718 734 72826 856
rect 72994 734 73102 856
rect 73270 734 73378 856
rect 73546 734 73654 856
rect 73822 734 73930 856
rect 74098 734 74206 856
rect 74374 734 74482 856
rect 74650 734 74758 856
rect 74926 734 75034 856
rect 75202 734 75310 856
rect 75478 734 75586 856
rect 75754 734 75862 856
rect 76030 734 76138 856
rect 76306 734 76414 856
rect 76582 734 76690 856
rect 76858 734 76966 856
rect 77134 734 77242 856
rect 77410 734 77518 856
rect 77686 734 77794 856
rect 77962 734 78070 856
rect 78238 734 78346 856
rect 78514 734 78622 856
rect 78790 734 78898 856
rect 79066 734 79174 856
rect 79342 734 79450 856
rect 79618 734 79726 856
rect 79894 734 80002 856
rect 80170 734 80278 856
rect 80446 734 80554 856
rect 80722 734 80830 856
rect 80998 734 81106 856
rect 81274 734 81382 856
rect 81550 734 81658 856
rect 81826 734 81934 856
rect 82102 734 82210 856
rect 82378 734 82486 856
rect 82654 734 82762 856
rect 82930 734 83038 856
rect 83206 734 83314 856
rect 83482 734 83590 856
rect 83758 734 83866 856
rect 84034 734 84142 856
rect 84310 734 84418 856
rect 84586 734 84694 856
rect 84862 734 84970 856
rect 85138 734 85246 856
rect 85414 734 85522 856
rect 85690 734 85798 856
rect 85966 734 86074 856
rect 86242 734 86350 856
rect 86518 734 86626 856
rect 86794 734 86902 856
rect 87070 734 87178 856
rect 87346 734 87454 856
rect 87622 734 87730 856
rect 87898 734 88006 856
rect 88174 734 88282 856
rect 88450 734 88558 856
rect 88726 734 88834 856
rect 89002 734 89110 856
rect 89278 734 89386 856
rect 89554 734 89662 856
rect 89830 734 89938 856
rect 90106 734 90214 856
rect 90382 734 90490 856
rect 90658 734 90766 856
rect 90934 734 91042 856
rect 91210 734 91318 856
rect 91486 734 91594 856
rect 91762 734 91870 856
rect 92038 734 92146 856
rect 92314 734 92422 856
rect 92590 734 92698 856
rect 92866 734 92974 856
rect 93142 734 93250 856
rect 93418 734 93526 856
rect 93694 734 93802 856
rect 93970 734 94078 856
rect 94246 734 94354 856
rect 94522 734 94630 856
rect 94798 734 94906 856
rect 95074 734 95182 856
rect 95350 734 95458 856
rect 95626 734 95734 856
rect 95902 734 96010 856
rect 96178 734 96286 856
rect 96454 734 96562 856
rect 96730 734 96838 856
rect 97006 734 97114 856
rect 97282 734 97390 856
rect 97558 734 97666 856
rect 97834 734 97942 856
rect 98110 734 98218 856
rect 98386 734 98494 856
rect 98662 734 98770 856
rect 98938 734 99046 856
rect 99214 734 99322 856
rect 99490 734 99598 856
rect 99766 734 99874 856
rect 100042 734 100150 856
rect 100318 734 100426 856
rect 100594 734 100702 856
rect 100870 734 100978 856
rect 101146 734 101254 856
rect 101422 734 101530 856
rect 101698 734 101806 856
rect 101974 734 102082 856
rect 102250 734 102358 856
rect 102526 734 102634 856
rect 102802 734 102910 856
rect 103078 734 103186 856
rect 103354 734 103462 856
rect 103630 734 103738 856
rect 103906 734 104014 856
rect 104182 734 104290 856
rect 104458 734 104566 856
rect 104734 734 104842 856
rect 105010 734 105118 856
rect 105286 734 105394 856
rect 105562 734 105670 856
rect 105838 734 105946 856
rect 106114 734 106222 856
rect 106390 734 106498 856
rect 106666 734 106774 856
rect 106942 734 107050 856
rect 107218 734 107326 856
rect 107494 734 107602 856
rect 107770 734 107878 856
rect 108046 734 108154 856
rect 108322 734 108430 856
rect 108598 734 108706 856
rect 108874 734 108982 856
rect 109150 734 109258 856
rect 109426 734 109534 856
rect 109702 734 109810 856
rect 109978 734 110086 856
rect 110254 734 110362 856
rect 110530 734 110638 856
rect 110806 734 110914 856
rect 111082 734 111190 856
rect 111358 734 111466 856
rect 111634 734 111742 856
rect 111910 734 112018 856
rect 112186 734 112294 856
rect 112462 734 112570 856
rect 112738 734 112846 856
rect 113014 734 113122 856
rect 113290 734 113398 856
rect 113566 734 113674 856
rect 113842 734 113950 856
rect 114118 734 114226 856
rect 114394 734 114502 856
rect 114670 734 114778 856
rect 114946 734 115054 856
rect 115222 734 115330 856
rect 115498 734 115606 856
rect 115774 734 115882 856
rect 116050 734 116158 856
rect 116326 734 116434 856
rect 116602 734 116710 856
rect 116878 734 116986 856
rect 117154 734 117262 856
rect 117430 734 117538 856
rect 117706 734 117814 856
rect 117982 734 118090 856
rect 118258 734 118366 856
rect 118534 734 118642 856
rect 118810 734 118918 856
rect 119086 734 119194 856
rect 119362 734 119470 856
rect 119638 734 119746 856
rect 119914 734 120022 856
rect 120190 734 120298 856
rect 120466 734 120574 856
rect 120742 734 120850 856
rect 121018 734 121126 856
rect 121294 734 121402 856
rect 121570 734 121678 856
rect 121846 734 121954 856
rect 122122 734 122230 856
rect 122398 734 122506 856
rect 122674 734 122782 856
rect 122950 734 123058 856
rect 123226 734 123334 856
rect 123502 734 123610 856
rect 123778 734 123886 856
rect 124054 734 124162 856
rect 124330 734 124438 856
rect 124606 734 124714 856
rect 124882 734 124990 856
rect 125158 734 125266 856
rect 125434 734 125542 856
rect 125710 734 125818 856
rect 125986 734 126094 856
rect 126262 734 126370 856
rect 126538 734 126646 856
rect 126814 734 126922 856
rect 127090 734 127198 856
rect 127366 734 127474 856
rect 127642 734 127750 856
rect 127918 734 128026 856
rect 128194 734 128302 856
rect 128470 734 128578 856
rect 128746 734 128854 856
rect 129022 734 129130 856
rect 129298 734 129406 856
rect 129574 734 129682 856
rect 129850 734 129958 856
rect 130126 734 130234 856
rect 130402 734 130510 856
rect 130678 734 130786 856
rect 130954 734 131062 856
rect 131230 734 131338 856
rect 131506 734 131614 856
rect 131782 734 131890 856
rect 132058 734 132166 856
rect 132334 734 132442 856
rect 132610 734 132718 856
rect 132886 734 132994 856
rect 133162 734 133270 856
rect 133438 734 133546 856
rect 133714 734 133822 856
rect 133990 734 134098 856
rect 134266 734 134374 856
rect 134542 734 134650 856
rect 134818 734 134926 856
rect 135094 734 135202 856
rect 135370 734 135478 856
rect 135646 734 135754 856
rect 135922 734 136030 856
rect 136198 734 136306 856
rect 136474 734 136582 856
rect 136750 734 136858 856
rect 137026 734 137134 856
rect 137302 734 137410 856
rect 137578 734 137686 856
rect 137854 734 137962 856
rect 138130 734 138238 856
rect 138406 734 138514 856
rect 138682 734 138790 856
rect 138958 734 139066 856
rect 139234 734 139342 856
rect 139510 734 139618 856
rect 139786 734 139894 856
rect 140062 734 140170 856
rect 140338 734 140446 856
rect 140614 734 140722 856
rect 140890 734 140998 856
rect 141166 734 141274 856
rect 141442 734 141550 856
rect 141718 734 141826 856
rect 141994 734 142102 856
rect 142270 734 142378 856
rect 142546 734 142654 856
rect 142822 734 142930 856
rect 143098 734 143206 856
rect 143374 734 143482 856
rect 143650 734 143758 856
rect 143926 734 144034 856
rect 144202 734 144310 856
rect 144478 734 144586 856
rect 144754 734 144862 856
rect 145030 734 145138 856
rect 145306 734 145414 856
rect 145582 734 145690 856
rect 145858 734 145966 856
rect 146134 734 146242 856
rect 146410 734 146518 856
rect 146686 734 146794 856
rect 146962 734 147070 856
rect 147238 734 147346 856
rect 147514 734 147622 856
rect 147790 734 147898 856
rect 148066 734 148174 856
rect 148342 734 148450 856
rect 148618 734 148726 856
rect 148894 734 149002 856
rect 149170 734 149278 856
rect 149446 734 149554 856
rect 149722 734 149830 856
rect 149998 734 150106 856
rect 150274 734 150382 856
rect 150550 734 150658 856
rect 150826 734 150934 856
rect 151102 734 151210 856
rect 151378 734 151486 856
rect 151654 734 151762 856
rect 151930 734 152038 856
rect 152206 734 152314 856
rect 152482 734 152590 856
rect 152758 734 152866 856
rect 153034 734 153142 856
rect 153310 734 153418 856
rect 153586 734 153694 856
rect 153862 734 153970 856
rect 154138 734 154246 856
rect 154414 734 154522 856
rect 154690 734 154798 856
rect 154966 734 155074 856
rect 155242 734 155350 856
rect 155518 734 155626 856
rect 155794 734 155902 856
rect 156070 734 156178 856
rect 156346 734 156454 856
rect 156622 734 156730 856
rect 156898 734 157006 856
rect 157174 734 157282 856
rect 157450 734 157558 856
rect 157726 734 157834 856
rect 158002 734 178314 856
<< obsm3 >>
rect 4210 2143 173486 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 1582 119200 1638 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48502 119200 48558 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 53194 119200 53250 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57886 119200 57942 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62578 119200 62634 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67270 119200 67326 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71962 119200 72018 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76654 119200 76710 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81346 119200 81402 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6274 119200 6330 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95422 119200 95478 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100114 119200 100170 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104806 119200 104862 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114190 119200 114246 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118882 119200 118938 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123574 119200 123630 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128266 119200 128322 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132958 119200 133014 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 137650 119200 137706 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10966 119200 11022 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142342 119200 142398 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147034 119200 147090 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 151726 119200 151782 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 156418 119200 156474 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161110 119200 161166 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165802 119200 165858 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 170494 119200 170550 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 175186 119200 175242 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 15658 119200 15714 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 20350 119200 20406 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 25042 119200 25098 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29734 119200 29790 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 34426 119200 34482 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 39118 119200 39174 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3146 119200 3202 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 50066 119200 50122 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54758 119200 54814 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68834 119200 68890 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73526 119200 73582 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78218 119200 78274 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82910 119200 82966 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101678 119200 101734 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111062 119200 111118 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115754 119200 115810 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120446 119200 120502 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125138 119200 125194 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129830 119200 129886 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134522 119200 134578 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139214 119200 139270 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143906 119200 143962 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 148598 119200 148654 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153290 119200 153346 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157982 119200 158038 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 162674 119200 162730 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172058 119200 172114 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176750 119200 176806 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21914 119200 21970 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26606 119200 26662 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 31298 119200 31354 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35990 119200 36046 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40682 119200 40738 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45374 119200 45430 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 119200 4766 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51630 119200 51686 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 56322 119200 56378 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 61014 119200 61070 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65706 119200 65762 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70398 119200 70454 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79782 119200 79838 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84474 119200 84530 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9402 119200 9458 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103242 119200 103298 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107934 119200 107990 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117318 119200 117374 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122010 119200 122066 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 126702 119200 126758 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131394 119200 131450 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140778 119200 140834 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 145470 119200 145526 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150162 119200 150218 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154854 119200 154910 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 159546 119200 159602 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168930 119200 168986 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 173622 119200 173678 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 178314 119200 178370 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18786 119200 18842 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 23478 119200 23534 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32862 119200 32918 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37554 119200 37610 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 42246 119200 42302 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 150990 0 151046 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 22098 0 22154 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7763560
string GDS_FILE /home/kareem_farid/cup_5-7-22/openlane/trainable_nn/runs/trainable_nn/results/signoff/trainable_nn.magic.gds
string GDS_START 391678
<< end >>

