magic
tech sky130A
magscale 1 2
timestamp 1670227627
<< nwell >>
rect 1066 156933 118902 157499
rect 1066 155845 118902 156411
rect 1066 154757 118902 155323
rect 1066 153669 118902 154235
rect 1066 152581 118902 153147
rect 1066 151493 118902 152059
rect 1066 150405 118902 150971
rect 1066 149317 118902 149883
rect 1066 148229 118902 148795
rect 1066 147141 118902 147707
rect 1066 146053 118902 146619
rect 1066 144965 118902 145531
rect 1066 143877 118902 144443
rect 1066 142789 118902 143355
rect 1066 141701 118902 142267
rect 1066 140613 118902 141179
rect 1066 139525 118902 140091
rect 1066 138437 118902 139003
rect 1066 137349 118902 137915
rect 1066 136261 118902 136827
rect 1066 135173 118902 135739
rect 1066 134085 118902 134651
rect 1066 132997 118902 133563
rect 1066 131909 118902 132475
rect 1066 130821 118902 131387
rect 1066 129733 118902 130299
rect 1066 128645 118902 129211
rect 1066 127557 118902 128123
rect 1066 126469 118902 127035
rect 1066 125381 118902 125947
rect 1066 124293 118902 124859
rect 1066 123205 118902 123771
rect 1066 122117 118902 122683
rect 1066 121029 118902 121595
rect 1066 119941 118902 120507
rect 1066 118853 118902 119419
rect 1066 117765 118902 118331
rect 1066 116677 118902 117243
rect 1066 115589 118902 116155
rect 1066 114501 118902 115067
rect 1066 113413 118902 113979
rect 1066 112325 118902 112891
rect 1066 111237 118902 111803
rect 1066 110149 118902 110715
rect 1066 109061 118902 109627
rect 1066 107973 118902 108539
rect 1066 106885 118902 107451
rect 1066 105797 118902 106363
rect 1066 104709 118902 105275
rect 1066 103621 118902 104187
rect 1066 102533 118902 103099
rect 1066 101445 118902 102011
rect 1066 100357 118902 100923
rect 1066 99269 118902 99835
rect 1066 98181 118902 98747
rect 1066 97093 118902 97659
rect 1066 96005 118902 96571
rect 1066 94917 118902 95483
rect 1066 93829 118902 94395
rect 1066 92741 118902 93307
rect 1066 91653 118902 92219
rect 1066 90565 118902 91131
rect 1066 89477 118902 90043
rect 1066 88389 118902 88955
rect 1066 87301 118902 87867
rect 1066 86213 118902 86779
rect 1066 85125 118902 85691
rect 1066 84037 118902 84603
rect 1066 82949 118902 83515
rect 1066 81861 118902 82427
rect 1066 80773 118902 81339
rect 1066 79685 118902 80251
rect 1066 78597 118902 79163
rect 1066 77509 118902 78075
rect 1066 76421 118902 76987
rect 1066 75333 118902 75899
rect 1066 74245 118902 74811
rect 1066 73157 118902 73723
rect 1066 72069 118902 72635
rect 1066 70981 118902 71547
rect 1066 69893 118902 70459
rect 1066 68805 118902 69371
rect 1066 67717 118902 68283
rect 1066 66629 118902 67195
rect 1066 65541 118902 66107
rect 1066 64453 118902 65019
rect 1066 63365 118902 63931
rect 1066 62277 118902 62843
rect 1066 61189 118902 61755
rect 1066 60101 118902 60667
rect 1066 59013 118902 59579
rect 1066 57925 118902 58491
rect 1066 56837 118902 57403
rect 1066 55749 118902 56315
rect 1066 54661 118902 55227
rect 1066 53573 118902 54139
rect 1066 52485 118902 53051
rect 1066 51397 118902 51963
rect 1066 50309 118902 50875
rect 1066 49221 118902 49787
rect 1066 48133 118902 48699
rect 1066 47045 118902 47611
rect 1066 45957 118902 46523
rect 1066 44869 118902 45435
rect 1066 43781 118902 44347
rect 1066 42693 118902 43259
rect 1066 41605 118902 42171
rect 1066 40517 118902 41083
rect 1066 39429 118902 39995
rect 1066 38341 118902 38907
rect 1066 37253 118902 37819
rect 1066 36165 118902 36731
rect 1066 35077 118902 35643
rect 1066 33989 118902 34555
rect 1066 32901 118902 33467
rect 1066 31813 118902 32379
rect 1066 30725 118902 31291
rect 1066 29637 118902 30203
rect 1066 28549 118902 29115
rect 1066 27461 118902 28027
rect 1066 26373 118902 26939
rect 1066 25285 118902 25851
rect 1066 24197 118902 24763
rect 1066 23109 118902 23675
rect 1066 22021 118902 22587
rect 1066 20933 118902 21499
rect 1066 19845 118902 20411
rect 1066 18757 118902 19323
rect 1066 17669 118902 18235
rect 1066 16581 118902 17147
rect 1066 15493 118902 16059
rect 1066 14405 118902 14971
rect 1066 13317 118902 13883
rect 1066 12229 118902 12795
rect 1066 11141 118902 11707
rect 1066 10053 118902 10619
rect 1066 8965 118902 9531
rect 1066 7877 118902 8443
rect 1066 6789 118902 7355
rect 1066 5701 118902 6267
rect 1066 4613 118902 5179
rect 1066 3525 118902 4091
rect 1066 2437 118902 3003
<< obsli1 >>
rect 1104 2159 118864 157777
<< obsm1 >>
rect 1104 8 119862 157808
<< metal2 >>
rect 2778 159200 2834 160000
rect 3790 159200 3846 160000
rect 4802 159200 4858 160000
rect 5814 159200 5870 160000
rect 6826 159200 6882 160000
rect 7838 159200 7894 160000
rect 8850 159200 8906 160000
rect 9862 159200 9918 160000
rect 10874 159200 10930 160000
rect 11886 159200 11942 160000
rect 12898 159200 12954 160000
rect 13910 159200 13966 160000
rect 14922 159200 14978 160000
rect 15934 159200 15990 160000
rect 16946 159200 17002 160000
rect 17958 159200 18014 160000
rect 18970 159200 19026 160000
rect 19982 159200 20038 160000
rect 20994 159200 21050 160000
rect 22006 159200 22062 160000
rect 23018 159200 23074 160000
rect 24030 159200 24086 160000
rect 25042 159200 25098 160000
rect 26054 159200 26110 160000
rect 27066 159200 27122 160000
rect 28078 159200 28134 160000
rect 29090 159200 29146 160000
rect 30102 159200 30158 160000
rect 31114 159200 31170 160000
rect 32126 159200 32182 160000
rect 33138 159200 33194 160000
rect 34150 159200 34206 160000
rect 35162 159200 35218 160000
rect 36174 159200 36230 160000
rect 37186 159200 37242 160000
rect 38198 159200 38254 160000
rect 39210 159200 39266 160000
rect 40222 159200 40278 160000
rect 41234 159200 41290 160000
rect 42246 159200 42302 160000
rect 43258 159200 43314 160000
rect 44270 159200 44326 160000
rect 45282 159200 45338 160000
rect 46294 159200 46350 160000
rect 47306 159200 47362 160000
rect 48318 159200 48374 160000
rect 49330 159200 49386 160000
rect 50342 159200 50398 160000
rect 51354 159200 51410 160000
rect 52366 159200 52422 160000
rect 53378 159200 53434 160000
rect 54390 159200 54446 160000
rect 55402 159200 55458 160000
rect 56414 159200 56470 160000
rect 57426 159200 57482 160000
rect 58438 159200 58494 160000
rect 59450 159200 59506 160000
rect 60462 159200 60518 160000
rect 61474 159200 61530 160000
rect 62486 159200 62542 160000
rect 63498 159200 63554 160000
rect 64510 159200 64566 160000
rect 65522 159200 65578 160000
rect 66534 159200 66590 160000
rect 67546 159200 67602 160000
rect 68558 159200 68614 160000
rect 69570 159200 69626 160000
rect 70582 159200 70638 160000
rect 71594 159200 71650 160000
rect 72606 159200 72662 160000
rect 73618 159200 73674 160000
rect 74630 159200 74686 160000
rect 75642 159200 75698 160000
rect 76654 159200 76710 160000
rect 77666 159200 77722 160000
rect 78678 159200 78734 160000
rect 79690 159200 79746 160000
rect 80702 159200 80758 160000
rect 81714 159200 81770 160000
rect 82726 159200 82782 160000
rect 83738 159200 83794 160000
rect 84750 159200 84806 160000
rect 85762 159200 85818 160000
rect 86774 159200 86830 160000
rect 87786 159200 87842 160000
rect 88798 159200 88854 160000
rect 89810 159200 89866 160000
rect 90822 159200 90878 160000
rect 91834 159200 91890 160000
rect 92846 159200 92902 160000
rect 93858 159200 93914 160000
rect 94870 159200 94926 160000
rect 95882 159200 95938 160000
rect 96894 159200 96950 160000
rect 97906 159200 97962 160000
rect 98918 159200 98974 160000
rect 99930 159200 99986 160000
rect 100942 159200 100998 160000
rect 101954 159200 102010 160000
rect 102966 159200 103022 160000
rect 103978 159200 104034 160000
rect 104990 159200 105046 160000
rect 106002 159200 106058 160000
rect 107014 159200 107070 160000
rect 108026 159200 108082 160000
rect 109038 159200 109094 160000
rect 110050 159200 110106 160000
rect 111062 159200 111118 160000
rect 112074 159200 112130 160000
rect 113086 159200 113142 160000
rect 114098 159200 114154 160000
rect 115110 159200 115166 160000
rect 116122 159200 116178 160000
rect 117134 159200 117190 160000
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98734 0 98790 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100022 0 100078 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102414 0 102470 800
rect 102598 0 102654 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104806 0 104862 800
rect 104990 0 105046 800
rect 105174 0 105230 800
<< obsm2 >>
rect 1306 159144 2722 159338
rect 2890 159144 3734 159338
rect 3902 159144 4746 159338
rect 4914 159144 5758 159338
rect 5926 159144 6770 159338
rect 6938 159144 7782 159338
rect 7950 159144 8794 159338
rect 8962 159144 9806 159338
rect 9974 159144 10818 159338
rect 10986 159144 11830 159338
rect 11998 159144 12842 159338
rect 13010 159144 13854 159338
rect 14022 159144 14866 159338
rect 15034 159144 15878 159338
rect 16046 159144 16890 159338
rect 17058 159144 17902 159338
rect 18070 159144 18914 159338
rect 19082 159144 19926 159338
rect 20094 159144 20938 159338
rect 21106 159144 21950 159338
rect 22118 159144 22962 159338
rect 23130 159144 23974 159338
rect 24142 159144 24986 159338
rect 25154 159144 25998 159338
rect 26166 159144 27010 159338
rect 27178 159144 28022 159338
rect 28190 159144 29034 159338
rect 29202 159144 30046 159338
rect 30214 159144 31058 159338
rect 31226 159144 32070 159338
rect 32238 159144 33082 159338
rect 33250 159144 34094 159338
rect 34262 159144 35106 159338
rect 35274 159144 36118 159338
rect 36286 159144 37130 159338
rect 37298 159144 38142 159338
rect 38310 159144 39154 159338
rect 39322 159144 40166 159338
rect 40334 159144 41178 159338
rect 41346 159144 42190 159338
rect 42358 159144 43202 159338
rect 43370 159144 44214 159338
rect 44382 159144 45226 159338
rect 45394 159144 46238 159338
rect 46406 159144 47250 159338
rect 47418 159144 48262 159338
rect 48430 159144 49274 159338
rect 49442 159144 50286 159338
rect 50454 159144 51298 159338
rect 51466 159144 52310 159338
rect 52478 159144 53322 159338
rect 53490 159144 54334 159338
rect 54502 159144 55346 159338
rect 55514 159144 56358 159338
rect 56526 159144 57370 159338
rect 57538 159144 58382 159338
rect 58550 159144 59394 159338
rect 59562 159144 60406 159338
rect 60574 159144 61418 159338
rect 61586 159144 62430 159338
rect 62598 159144 63442 159338
rect 63610 159144 64454 159338
rect 64622 159144 65466 159338
rect 65634 159144 66478 159338
rect 66646 159144 67490 159338
rect 67658 159144 68502 159338
rect 68670 159144 69514 159338
rect 69682 159144 70526 159338
rect 70694 159144 71538 159338
rect 71706 159144 72550 159338
rect 72718 159144 73562 159338
rect 73730 159144 74574 159338
rect 74742 159144 75586 159338
rect 75754 159144 76598 159338
rect 76766 159144 77610 159338
rect 77778 159144 78622 159338
rect 78790 159144 79634 159338
rect 79802 159144 80646 159338
rect 80814 159144 81658 159338
rect 81826 159144 82670 159338
rect 82838 159144 83682 159338
rect 83850 159144 84694 159338
rect 84862 159144 85706 159338
rect 85874 159144 86718 159338
rect 86886 159144 87730 159338
rect 87898 159144 88742 159338
rect 88910 159144 89754 159338
rect 89922 159144 90766 159338
rect 90934 159144 91778 159338
rect 91946 159144 92790 159338
rect 92958 159144 93802 159338
rect 93970 159144 94814 159338
rect 94982 159144 95826 159338
rect 95994 159144 96838 159338
rect 97006 159144 97850 159338
rect 98018 159144 98862 159338
rect 99030 159144 99874 159338
rect 100042 159144 100886 159338
rect 101054 159144 101898 159338
rect 102066 159144 102910 159338
rect 103078 159144 103922 159338
rect 104090 159144 104934 159338
rect 105102 159144 105946 159338
rect 106114 159144 106958 159338
rect 107126 159144 107970 159338
rect 108138 159144 108982 159338
rect 109150 159144 109994 159338
rect 110162 159144 111006 159338
rect 111174 159144 112018 159338
rect 112186 159144 113030 159338
rect 113198 159144 114042 159338
rect 114210 159144 115054 159338
rect 115222 159144 116066 159338
rect 116234 159144 117078 159338
rect 117246 159144 119856 159338
rect 1306 856 119856 159144
rect 1306 2 14590 856
rect 14758 2 14774 856
rect 14942 2 14958 856
rect 15126 2 15142 856
rect 15310 2 15326 856
rect 15494 2 15510 856
rect 15678 2 15694 856
rect 15862 2 15878 856
rect 16046 2 16062 856
rect 16230 2 16246 856
rect 16414 2 16430 856
rect 16598 2 16614 856
rect 16782 2 16798 856
rect 16966 2 16982 856
rect 17150 2 17166 856
rect 17334 2 17350 856
rect 17518 2 17534 856
rect 17702 2 17718 856
rect 17886 2 17902 856
rect 18070 2 18086 856
rect 18254 2 18270 856
rect 18438 2 18454 856
rect 18622 2 18638 856
rect 18806 2 18822 856
rect 18990 2 19006 856
rect 19174 2 19190 856
rect 19358 2 19374 856
rect 19542 2 19558 856
rect 19726 2 19742 856
rect 19910 2 19926 856
rect 20094 2 20110 856
rect 20278 2 20294 856
rect 20462 2 20478 856
rect 20646 2 20662 856
rect 20830 2 20846 856
rect 21014 2 21030 856
rect 21198 2 21214 856
rect 21382 2 21398 856
rect 21566 2 21582 856
rect 21750 2 21766 856
rect 21934 2 21950 856
rect 22118 2 22134 856
rect 22302 2 22318 856
rect 22486 2 22502 856
rect 22670 2 22686 856
rect 22854 2 22870 856
rect 23038 2 23054 856
rect 23222 2 23238 856
rect 23406 2 23422 856
rect 23590 2 23606 856
rect 23774 2 23790 856
rect 23958 2 23974 856
rect 24142 2 24158 856
rect 24326 2 24342 856
rect 24510 2 24526 856
rect 24694 2 24710 856
rect 24878 2 24894 856
rect 25062 2 25078 856
rect 25246 2 25262 856
rect 25430 2 25446 856
rect 25614 2 25630 856
rect 25798 2 25814 856
rect 25982 2 25998 856
rect 26166 2 26182 856
rect 26350 2 26366 856
rect 26534 2 26550 856
rect 26718 2 26734 856
rect 26902 2 26918 856
rect 27086 2 27102 856
rect 27270 2 27286 856
rect 27454 2 27470 856
rect 27638 2 27654 856
rect 27822 2 27838 856
rect 28006 2 28022 856
rect 28190 2 28206 856
rect 28374 2 28390 856
rect 28558 2 28574 856
rect 28742 2 28758 856
rect 28926 2 28942 856
rect 29110 2 29126 856
rect 29294 2 29310 856
rect 29478 2 29494 856
rect 29662 2 29678 856
rect 29846 2 29862 856
rect 30030 2 30046 856
rect 30214 2 30230 856
rect 30398 2 30414 856
rect 30582 2 30598 856
rect 30766 2 30782 856
rect 30950 2 30966 856
rect 31134 2 31150 856
rect 31318 2 31334 856
rect 31502 2 31518 856
rect 31686 2 31702 856
rect 31870 2 31886 856
rect 32054 2 32070 856
rect 32238 2 32254 856
rect 32422 2 32438 856
rect 32606 2 32622 856
rect 32790 2 32806 856
rect 32974 2 32990 856
rect 33158 2 33174 856
rect 33342 2 33358 856
rect 33526 2 33542 856
rect 33710 2 33726 856
rect 33894 2 33910 856
rect 34078 2 34094 856
rect 34262 2 34278 856
rect 34446 2 34462 856
rect 34630 2 34646 856
rect 34814 2 34830 856
rect 34998 2 35014 856
rect 35182 2 35198 856
rect 35366 2 35382 856
rect 35550 2 35566 856
rect 35734 2 35750 856
rect 35918 2 35934 856
rect 36102 2 36118 856
rect 36286 2 36302 856
rect 36470 2 36486 856
rect 36654 2 36670 856
rect 36838 2 36854 856
rect 37022 2 37038 856
rect 37206 2 37222 856
rect 37390 2 37406 856
rect 37574 2 37590 856
rect 37758 2 37774 856
rect 37942 2 37958 856
rect 38126 2 38142 856
rect 38310 2 38326 856
rect 38494 2 38510 856
rect 38678 2 38694 856
rect 38862 2 38878 856
rect 39046 2 39062 856
rect 39230 2 39246 856
rect 39414 2 39430 856
rect 39598 2 39614 856
rect 39782 2 39798 856
rect 39966 2 39982 856
rect 40150 2 40166 856
rect 40334 2 40350 856
rect 40518 2 40534 856
rect 40702 2 40718 856
rect 40886 2 40902 856
rect 41070 2 41086 856
rect 41254 2 41270 856
rect 41438 2 41454 856
rect 41622 2 41638 856
rect 41806 2 41822 856
rect 41990 2 42006 856
rect 42174 2 42190 856
rect 42358 2 42374 856
rect 42542 2 42558 856
rect 42726 2 42742 856
rect 42910 2 42926 856
rect 43094 2 43110 856
rect 43278 2 43294 856
rect 43462 2 43478 856
rect 43646 2 43662 856
rect 43830 2 43846 856
rect 44014 2 44030 856
rect 44198 2 44214 856
rect 44382 2 44398 856
rect 44566 2 44582 856
rect 44750 2 44766 856
rect 44934 2 44950 856
rect 45118 2 45134 856
rect 45302 2 45318 856
rect 45486 2 45502 856
rect 45670 2 45686 856
rect 45854 2 45870 856
rect 46038 2 46054 856
rect 46222 2 46238 856
rect 46406 2 46422 856
rect 46590 2 46606 856
rect 46774 2 46790 856
rect 46958 2 46974 856
rect 47142 2 47158 856
rect 47326 2 47342 856
rect 47510 2 47526 856
rect 47694 2 47710 856
rect 47878 2 47894 856
rect 48062 2 48078 856
rect 48246 2 48262 856
rect 48430 2 48446 856
rect 48614 2 48630 856
rect 48798 2 48814 856
rect 48982 2 48998 856
rect 49166 2 49182 856
rect 49350 2 49366 856
rect 49534 2 49550 856
rect 49718 2 49734 856
rect 49902 2 49918 856
rect 50086 2 50102 856
rect 50270 2 50286 856
rect 50454 2 50470 856
rect 50638 2 50654 856
rect 50822 2 50838 856
rect 51006 2 51022 856
rect 51190 2 51206 856
rect 51374 2 51390 856
rect 51558 2 51574 856
rect 51742 2 51758 856
rect 51926 2 51942 856
rect 52110 2 52126 856
rect 52294 2 52310 856
rect 52478 2 52494 856
rect 52662 2 52678 856
rect 52846 2 52862 856
rect 53030 2 53046 856
rect 53214 2 53230 856
rect 53398 2 53414 856
rect 53582 2 53598 856
rect 53766 2 53782 856
rect 53950 2 53966 856
rect 54134 2 54150 856
rect 54318 2 54334 856
rect 54502 2 54518 856
rect 54686 2 54702 856
rect 54870 2 54886 856
rect 55054 2 55070 856
rect 55238 2 55254 856
rect 55422 2 55438 856
rect 55606 2 55622 856
rect 55790 2 55806 856
rect 55974 2 55990 856
rect 56158 2 56174 856
rect 56342 2 56358 856
rect 56526 2 56542 856
rect 56710 2 56726 856
rect 56894 2 56910 856
rect 57078 2 57094 856
rect 57262 2 57278 856
rect 57446 2 57462 856
rect 57630 2 57646 856
rect 57814 2 57830 856
rect 57998 2 58014 856
rect 58182 2 58198 856
rect 58366 2 58382 856
rect 58550 2 58566 856
rect 58734 2 58750 856
rect 58918 2 58934 856
rect 59102 2 59118 856
rect 59286 2 59302 856
rect 59470 2 59486 856
rect 59654 2 59670 856
rect 59838 2 59854 856
rect 60022 2 60038 856
rect 60206 2 60222 856
rect 60390 2 60406 856
rect 60574 2 60590 856
rect 60758 2 60774 856
rect 60942 2 60958 856
rect 61126 2 61142 856
rect 61310 2 61326 856
rect 61494 2 61510 856
rect 61678 2 61694 856
rect 61862 2 61878 856
rect 62046 2 62062 856
rect 62230 2 62246 856
rect 62414 2 62430 856
rect 62598 2 62614 856
rect 62782 2 62798 856
rect 62966 2 62982 856
rect 63150 2 63166 856
rect 63334 2 63350 856
rect 63518 2 63534 856
rect 63702 2 63718 856
rect 63886 2 63902 856
rect 64070 2 64086 856
rect 64254 2 64270 856
rect 64438 2 64454 856
rect 64622 2 64638 856
rect 64806 2 64822 856
rect 64990 2 65006 856
rect 65174 2 65190 856
rect 65358 2 65374 856
rect 65542 2 65558 856
rect 65726 2 65742 856
rect 65910 2 65926 856
rect 66094 2 66110 856
rect 66278 2 66294 856
rect 66462 2 66478 856
rect 66646 2 66662 856
rect 66830 2 66846 856
rect 67014 2 67030 856
rect 67198 2 67214 856
rect 67382 2 67398 856
rect 67566 2 67582 856
rect 67750 2 67766 856
rect 67934 2 67950 856
rect 68118 2 68134 856
rect 68302 2 68318 856
rect 68486 2 68502 856
rect 68670 2 68686 856
rect 68854 2 68870 856
rect 69038 2 69054 856
rect 69222 2 69238 856
rect 69406 2 69422 856
rect 69590 2 69606 856
rect 69774 2 69790 856
rect 69958 2 69974 856
rect 70142 2 70158 856
rect 70326 2 70342 856
rect 70510 2 70526 856
rect 70694 2 70710 856
rect 70878 2 70894 856
rect 71062 2 71078 856
rect 71246 2 71262 856
rect 71430 2 71446 856
rect 71614 2 71630 856
rect 71798 2 71814 856
rect 71982 2 71998 856
rect 72166 2 72182 856
rect 72350 2 72366 856
rect 72534 2 72550 856
rect 72718 2 72734 856
rect 72902 2 72918 856
rect 73086 2 73102 856
rect 73270 2 73286 856
rect 73454 2 73470 856
rect 73638 2 73654 856
rect 73822 2 73838 856
rect 74006 2 74022 856
rect 74190 2 74206 856
rect 74374 2 74390 856
rect 74558 2 74574 856
rect 74742 2 74758 856
rect 74926 2 74942 856
rect 75110 2 75126 856
rect 75294 2 75310 856
rect 75478 2 75494 856
rect 75662 2 75678 856
rect 75846 2 75862 856
rect 76030 2 76046 856
rect 76214 2 76230 856
rect 76398 2 76414 856
rect 76582 2 76598 856
rect 76766 2 76782 856
rect 76950 2 76966 856
rect 77134 2 77150 856
rect 77318 2 77334 856
rect 77502 2 77518 856
rect 77686 2 77702 856
rect 77870 2 77886 856
rect 78054 2 78070 856
rect 78238 2 78254 856
rect 78422 2 78438 856
rect 78606 2 78622 856
rect 78790 2 78806 856
rect 78974 2 78990 856
rect 79158 2 79174 856
rect 79342 2 79358 856
rect 79526 2 79542 856
rect 79710 2 79726 856
rect 79894 2 79910 856
rect 80078 2 80094 856
rect 80262 2 80278 856
rect 80446 2 80462 856
rect 80630 2 80646 856
rect 80814 2 80830 856
rect 80998 2 81014 856
rect 81182 2 81198 856
rect 81366 2 81382 856
rect 81550 2 81566 856
rect 81734 2 81750 856
rect 81918 2 81934 856
rect 82102 2 82118 856
rect 82286 2 82302 856
rect 82470 2 82486 856
rect 82654 2 82670 856
rect 82838 2 82854 856
rect 83022 2 83038 856
rect 83206 2 83222 856
rect 83390 2 83406 856
rect 83574 2 83590 856
rect 83758 2 83774 856
rect 83942 2 83958 856
rect 84126 2 84142 856
rect 84310 2 84326 856
rect 84494 2 84510 856
rect 84678 2 84694 856
rect 84862 2 84878 856
rect 85046 2 85062 856
rect 85230 2 85246 856
rect 85414 2 85430 856
rect 85598 2 85614 856
rect 85782 2 85798 856
rect 85966 2 85982 856
rect 86150 2 86166 856
rect 86334 2 86350 856
rect 86518 2 86534 856
rect 86702 2 86718 856
rect 86886 2 86902 856
rect 87070 2 87086 856
rect 87254 2 87270 856
rect 87438 2 87454 856
rect 87622 2 87638 856
rect 87806 2 87822 856
rect 87990 2 88006 856
rect 88174 2 88190 856
rect 88358 2 88374 856
rect 88542 2 88558 856
rect 88726 2 88742 856
rect 88910 2 88926 856
rect 89094 2 89110 856
rect 89278 2 89294 856
rect 89462 2 89478 856
rect 89646 2 89662 856
rect 89830 2 89846 856
rect 90014 2 90030 856
rect 90198 2 90214 856
rect 90382 2 90398 856
rect 90566 2 90582 856
rect 90750 2 90766 856
rect 90934 2 90950 856
rect 91118 2 91134 856
rect 91302 2 91318 856
rect 91486 2 91502 856
rect 91670 2 91686 856
rect 91854 2 91870 856
rect 92038 2 92054 856
rect 92222 2 92238 856
rect 92406 2 92422 856
rect 92590 2 92606 856
rect 92774 2 92790 856
rect 92958 2 92974 856
rect 93142 2 93158 856
rect 93326 2 93342 856
rect 93510 2 93526 856
rect 93694 2 93710 856
rect 93878 2 93894 856
rect 94062 2 94078 856
rect 94246 2 94262 856
rect 94430 2 94446 856
rect 94614 2 94630 856
rect 94798 2 94814 856
rect 94982 2 94998 856
rect 95166 2 95182 856
rect 95350 2 95366 856
rect 95534 2 95550 856
rect 95718 2 95734 856
rect 95902 2 95918 856
rect 96086 2 96102 856
rect 96270 2 96286 856
rect 96454 2 96470 856
rect 96638 2 96654 856
rect 96822 2 96838 856
rect 97006 2 97022 856
rect 97190 2 97206 856
rect 97374 2 97390 856
rect 97558 2 97574 856
rect 97742 2 97758 856
rect 97926 2 97942 856
rect 98110 2 98126 856
rect 98294 2 98310 856
rect 98478 2 98494 856
rect 98662 2 98678 856
rect 98846 2 98862 856
rect 99030 2 99046 856
rect 99214 2 99230 856
rect 99398 2 99414 856
rect 99582 2 99598 856
rect 99766 2 99782 856
rect 99950 2 99966 856
rect 100134 2 100150 856
rect 100318 2 100334 856
rect 100502 2 100518 856
rect 100686 2 100702 856
rect 100870 2 100886 856
rect 101054 2 101070 856
rect 101238 2 101254 856
rect 101422 2 101438 856
rect 101606 2 101622 856
rect 101790 2 101806 856
rect 101974 2 101990 856
rect 102158 2 102174 856
rect 102342 2 102358 856
rect 102526 2 102542 856
rect 102710 2 102726 856
rect 102894 2 102910 856
rect 103078 2 103094 856
rect 103262 2 103278 856
rect 103446 2 103462 856
rect 103630 2 103646 856
rect 103814 2 103830 856
rect 103998 2 104014 856
rect 104182 2 104198 856
rect 104366 2 104382 856
rect 104550 2 104566 856
rect 104734 2 104750 856
rect 104918 2 104934 856
rect 105102 2 105118 856
rect 105286 2 119856 856
<< obsm3 >>
rect 1301 443 119495 157793
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< obsm4 >>
rect 1715 2048 4128 153509
rect 4608 2048 19488 153509
rect 19968 2048 34848 153509
rect 35328 2048 50208 153509
rect 50688 2048 65568 153509
rect 66048 2048 80928 153509
rect 81408 2048 96288 153509
rect 96768 2048 111648 153509
rect 112128 2048 117333 153509
rect 1715 443 117333 2048
<< labels >>
rlabel metal2 s 2778 159200 2834 160000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 33138 159200 33194 160000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 36174 159200 36230 160000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 39210 159200 39266 160000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 42246 159200 42302 160000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 45282 159200 45338 160000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 48318 159200 48374 160000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 51354 159200 51410 160000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 54390 159200 54446 160000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 57426 159200 57482 160000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 60462 159200 60518 160000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5814 159200 5870 160000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 63498 159200 63554 160000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 66534 159200 66590 160000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 69570 159200 69626 160000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 72606 159200 72662 160000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 75642 159200 75698 160000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 78678 159200 78734 160000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 81714 159200 81770 160000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 84750 159200 84806 160000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 87786 159200 87842 160000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 90822 159200 90878 160000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 8850 159200 8906 160000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 93858 159200 93914 160000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 96894 159200 96950 160000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 99930 159200 99986 160000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 102966 159200 103022 160000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 106002 159200 106058 160000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 109038 159200 109094 160000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 112074 159200 112130 160000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 115110 159200 115166 160000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 11886 159200 11942 160000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 14922 159200 14978 160000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 17958 159200 18014 160000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 20994 159200 21050 160000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 24030 159200 24086 160000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 27066 159200 27122 160000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 30102 159200 30158 160000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3790 159200 3846 160000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 34150 159200 34206 160000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 37186 159200 37242 160000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 40222 159200 40278 160000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 43258 159200 43314 160000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 46294 159200 46350 160000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 49330 159200 49386 160000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 52366 159200 52422 160000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 55402 159200 55458 160000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 58438 159200 58494 160000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 61474 159200 61530 160000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6826 159200 6882 160000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 64510 159200 64566 160000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 67546 159200 67602 160000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70582 159200 70638 160000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 73618 159200 73674 160000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 76654 159200 76710 160000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 79690 159200 79746 160000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 82726 159200 82782 160000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 85762 159200 85818 160000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 88798 159200 88854 160000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 91834 159200 91890 160000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 9862 159200 9918 160000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 94870 159200 94926 160000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 97906 159200 97962 160000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 100942 159200 100998 160000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 103978 159200 104034 160000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 107014 159200 107070 160000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 110050 159200 110106 160000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 113086 159200 113142 160000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 116122 159200 116178 160000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 12898 159200 12954 160000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 15934 159200 15990 160000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 18970 159200 19026 160000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 22006 159200 22062 160000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 25042 159200 25098 160000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 28078 159200 28134 160000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 31114 159200 31170 160000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4802 159200 4858 160000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 35162 159200 35218 160000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 38198 159200 38254 160000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 41234 159200 41290 160000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 44270 159200 44326 160000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 47306 159200 47362 160000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 50342 159200 50398 160000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 53378 159200 53434 160000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 56414 159200 56470 160000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 59450 159200 59506 160000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 62486 159200 62542 160000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7838 159200 7894 160000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 65522 159200 65578 160000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 68558 159200 68614 160000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 71594 159200 71650 160000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 74630 159200 74686 160000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 77666 159200 77722 160000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 80702 159200 80758 160000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 83738 159200 83794 160000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 86774 159200 86830 160000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 89810 159200 89866 160000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 92846 159200 92902 160000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 10874 159200 10930 160000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 95882 159200 95938 160000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 98918 159200 98974 160000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 101954 159200 102010 160000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 104990 159200 105046 160000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 108026 159200 108082 160000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 111062 159200 111118 160000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 114098 159200 114154 160000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 117134 159200 117190 160000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 13910 159200 13966 160000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 16946 159200 17002 160000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 19982 159200 20038 160000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 23018 159200 23074 160000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 26054 159200 26110 160000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 29090 159200 29146 160000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 32126 159200 32182 160000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 105174 0 105230 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 14646 0 14702 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 60199312
string GDS_FILE /home/htamas/progs/trainable-nn-resub2/openlane/trainable_nn/runs/22_12_05_08_19/results/signoff/trainable_nn.magic.gds
string GDS_START 1396014
<< end >>

