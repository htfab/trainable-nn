magic
tech sky130B
magscale 1 2
timestamp 1663048546
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 283834 700884 283840 700936
rect 283892 700924 283898 700936
rect 301406 700924 301412 700936
rect 283892 700896 301412 700924
rect 283892 700884 283898 700896
rect 301406 700884 301412 700896
rect 301464 700884 301470 700936
rect 290090 700816 290096 700868
rect 290148 700856 290154 700868
rect 348786 700856 348792 700868
rect 290148 700828 348792 700856
rect 290148 700816 290154 700828
rect 348786 700816 348792 700828
rect 348844 700816 348850 700868
rect 218974 700748 218980 700800
rect 219032 700788 219038 700800
rect 312722 700788 312728 700800
rect 219032 700760 312728 700788
rect 219032 700748 219038 700760
rect 312722 700748 312728 700760
rect 312780 700748 312786 700800
rect 278774 700680 278780 700732
rect 278832 700720 278838 700732
rect 413646 700720 413652 700732
rect 278832 700692 413652 700720
rect 278832 700680 278838 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 324038 700652 324044 700664
rect 154172 700624 324044 700652
rect 154172 700612 154178 700624
rect 324038 700612 324044 700624
rect 324096 700612 324102 700664
rect 267458 700544 267464 700596
rect 267516 700584 267522 700596
rect 478506 700584 478512 700596
rect 267516 700556 478512 700584
rect 267516 700544 267522 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 335354 700516 335360 700528
rect 89220 700488 335360 700516
rect 89220 700476 89226 700488
rect 335354 700476 335360 700488
rect 335412 700476 335418 700528
rect 256142 700408 256148 700460
rect 256200 700448 256206 700460
rect 543458 700448 543464 700460
rect 256200 700420 543464 700448
rect 256200 700408 256206 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 346670 700380 346676 700392
rect 24360 700352 346676 700380
rect 24360 700340 24366 700352
rect 346670 700340 346676 700352
rect 346728 700340 346734 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 342898 700312 342904 700324
rect 8168 700284 342904 700312
rect 8168 700272 8174 700284
rect 342898 700272 342904 700284
rect 342956 700272 342962 700324
rect 549898 700272 549904 700324
rect 549956 700312 549962 700324
rect 559650 700312 559656 700324
rect 549956 700284 559656 700312
rect 549956 700272 549962 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 267642 698980 267648 699032
rect 267700 699020 267706 699032
rect 297634 699020 297640 699032
rect 267700 698992 297640 699020
rect 267700 698980 267706 698992
rect 297634 698980 297640 698992
rect 297692 698980 297698 699032
rect 275002 698912 275008 698964
rect 275060 698952 275066 698964
rect 397454 698952 397460 698964
rect 275060 698924 397460 698952
rect 275060 698912 275066 698924
rect 397454 698912 397460 698924
rect 397512 698912 397518 698964
rect 137830 697552 137836 697604
rect 137888 697592 137894 697604
rect 320266 697592 320272 697604
rect 137888 697564 320272 697592
rect 137888 697552 137894 697564
rect 320266 697552 320272 697564
rect 320324 697552 320330 697604
rect 241054 696940 241060 696992
rect 241112 696980 241118 696992
rect 580166 696980 580172 696992
rect 241112 696952 580172 696980
rect 241112 696940 241118 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 105446 696192 105452 696244
rect 105504 696232 105510 696244
rect 327810 696232 327816 696244
rect 105504 696204 327816 696232
rect 105504 696192 105510 696204
rect 327810 696192 327816 696204
rect 327868 696192 327874 696244
rect 244826 683204 244832 683256
rect 244884 683244 244890 683256
rect 580166 683244 580172 683256
rect 244884 683216 580172 683244
rect 244884 683204 244890 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 350442 683176 350448 683188
rect 3476 683148 350448 683176
rect 3476 683136 3482 683148
rect 350442 683136 350448 683148
rect 350500 683136 350506 683188
rect 237282 670760 237288 670812
rect 237340 670800 237346 670812
rect 580166 670800 580172 670812
rect 237340 670772 580172 670800
rect 237340 670760 237346 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 357986 670732 357992 670744
rect 3568 670704 357992 670732
rect 3568 670692 3574 670704
rect 357986 670692 357992 670704
rect 358044 670692 358050 670744
rect 286318 663008 286324 663060
rect 286376 663048 286382 663060
rect 331214 663048 331220 663060
rect 286376 663020 331220 663048
rect 286376 663008 286382 663020
rect 331214 663008 331220 663020
rect 331272 663008 331278 663060
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 354214 656928 354220 656940
rect 3476 656900 354220 656928
rect 3476 656888 3482 656900
rect 354214 656888 354220 656900
rect 354272 656888 354278 656940
rect 229738 643084 229744 643136
rect 229796 643124 229802 643136
rect 580166 643124 580172 643136
rect 229796 643096 580172 643124
rect 229796 643084 229802 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 201494 642336 201500 642388
rect 201552 642376 201558 642388
rect 308950 642376 308956 642388
rect 201552 642348 308956 642376
rect 201552 642336 201558 642348
rect 308950 642336 308956 642348
rect 309008 642336 309014 642388
rect 234614 640976 234620 641028
rect 234672 641016 234678 641028
rect 305178 641016 305184 641028
rect 234672 640988 305184 641016
rect 234672 640976 234678 640988
rect 305178 640976 305184 640988
rect 305236 640976 305242 641028
rect 263686 639548 263692 639600
rect 263744 639588 263750 639600
rect 462314 639588 462320 639600
rect 263744 639560 462320 639588
rect 263744 639548 263750 639560
rect 462314 639548 462320 639560
rect 462372 639548 462378 639600
rect 71774 638392 71780 638444
rect 71832 638432 71838 638444
rect 331582 638432 331588 638444
rect 71832 638404 331588 638432
rect 71832 638392 71838 638404
rect 331582 638392 331588 638404
rect 331640 638392 331646 638444
rect 252370 638324 252376 638376
rect 252428 638364 252434 638376
rect 527174 638364 527180 638376
rect 252428 638336 527180 638364
rect 252428 638324 252434 638336
rect 527174 638324 527180 638336
rect 527232 638324 527238 638376
rect 68370 638256 68376 638308
rect 68428 638296 68434 638308
rect 369302 638296 369308 638308
rect 68428 638268 369308 638296
rect 68428 638256 68434 638268
rect 369302 638256 369308 638268
rect 369360 638256 369366 638308
rect 184474 638188 184480 638240
rect 184532 638228 184538 638240
rect 522390 638228 522396 638240
rect 184532 638200 522396 638228
rect 184532 638188 184538 638200
rect 522390 638188 522396 638200
rect 522448 638188 522454 638240
rect 58618 638120 58624 638172
rect 58676 638160 58682 638172
rect 403250 638160 403256 638172
rect 58676 638132 403256 638160
rect 58676 638120 58682 638132
rect 403250 638120 403256 638132
rect 403308 638120 403314 638172
rect 173158 638052 173164 638104
rect 173216 638092 173222 638104
rect 521010 638092 521016 638104
rect 173216 638064 521016 638092
rect 173216 638052 173222 638064
rect 521010 638052 521016 638064
rect 521068 638052 521074 638104
rect 161842 637984 161848 638036
rect 161900 638024 161906 638036
rect 520918 638024 520924 638036
rect 161900 637996 520924 638024
rect 161900 637984 161906 637996
rect 520918 637984 520924 637996
rect 520976 637984 520982 638036
rect 57238 637916 57244 637968
rect 57296 637956 57302 637968
rect 422110 637956 422116 637968
rect 57296 637928 422116 637956
rect 57296 637916 57302 637928
rect 422110 637916 422116 637928
rect 422168 637916 422174 637968
rect 150526 637848 150532 637900
rect 150584 637888 150590 637900
rect 518250 637888 518256 637900
rect 150584 637860 518256 637888
rect 150584 637848 150590 637860
rect 518250 637848 518256 637860
rect 518308 637848 518314 637900
rect 7558 637780 7564 637832
rect 7616 637820 7622 637832
rect 388162 637820 388168 637832
rect 7616 637792 388168 637820
rect 7616 637780 7622 637792
rect 388162 637780 388168 637792
rect 388220 637780 388226 637832
rect 13078 637712 13084 637764
rect 13136 637752 13142 637764
rect 410426 637752 410432 637764
rect 13136 637724 410432 637752
rect 13136 637712 13142 637724
rect 410426 637712 410432 637724
rect 410484 637712 410490 637764
rect 109034 637644 109040 637696
rect 109092 637684 109098 637696
rect 515398 637684 515404 637696
rect 109092 637656 515404 637684
rect 109092 637644 109098 637656
rect 515398 637644 515404 637656
rect 515456 637644 515462 637696
rect 105262 637576 105268 637628
rect 105320 637616 105326 637628
rect 516778 637616 516784 637628
rect 105320 637588 516784 637616
rect 105320 637576 105326 637588
rect 516778 637576 516784 637588
rect 516836 637576 516842 637628
rect 169754 637100 169760 637152
rect 169812 637140 169818 637152
rect 316126 637140 316132 637152
rect 169812 637112 316132 637140
rect 169812 637100 169818 637112
rect 316126 637100 316132 637112
rect 316184 637100 316190 637152
rect 40034 637032 40040 637084
rect 40092 637072 40098 637084
rect 338758 637072 338764 637084
rect 40092 637044 338764 637072
rect 40092 637032 40098 637044
rect 338758 637032 338764 637044
rect 338816 637032 338822 637084
rect 248874 636964 248880 637016
rect 248932 637004 248938 637016
rect 549898 637004 549904 637016
rect 248932 636976 549904 637004
rect 248932 636964 248938 636976
rect 549898 636964 549904 636976
rect 549956 636964 549962 637016
rect 180702 636896 180708 636948
rect 180760 636936 180766 636948
rect 516962 636936 516968 636948
rect 180760 636908 516968 636936
rect 180760 636896 180766 636908
rect 516962 636896 516968 636908
rect 517020 636896 517026 636948
rect 53098 636828 53104 636880
rect 53156 636868 53162 636880
rect 414198 636868 414204 636880
rect 53156 636840 414204 636868
rect 53156 636828 53162 636840
rect 414198 636828 414204 636840
rect 414256 636828 414262 636880
rect 147030 636760 147036 636812
rect 147088 636800 147094 636812
rect 516870 636800 516876 636812
rect 147088 636772 516876 636800
rect 147088 636760 147094 636772
rect 516870 636760 516876 636772
rect 516928 636760 516934 636812
rect 66898 636692 66904 636744
rect 66956 636732 66962 636744
rect 440602 636732 440608 636744
rect 66956 636704 440608 636732
rect 66956 636692 66962 636704
rect 440602 636692 440608 636704
rect 440660 636692 440666 636744
rect 124122 636624 124128 636676
rect 124180 636664 124186 636676
rect 514202 636664 514208 636676
rect 124180 636636 514208 636664
rect 124180 636624 124186 636636
rect 514202 636624 514208 636636
rect 514260 636624 514266 636676
rect 71038 636556 71044 636608
rect 71096 636596 71102 636608
rect 463234 636596 463240 636608
rect 71096 636568 463240 636596
rect 71096 636556 71102 636568
rect 463234 636556 463240 636568
rect 463292 636556 463298 636608
rect 64138 636488 64144 636540
rect 64196 636528 64202 636540
rect 474734 636528 474740 636540
rect 64196 636500 474740 636528
rect 64196 636488 64202 636500
rect 474734 636488 474740 636500
rect 474792 636488 474798 636540
rect 68278 636420 68284 636472
rect 68336 636460 68342 636472
rect 485866 636460 485872 636472
rect 68336 636432 485872 636460
rect 68336 636420 68342 636432
rect 485866 636420 485872 636432
rect 485924 636420 485930 636472
rect 72418 636352 72424 636404
rect 72476 636392 72482 636404
rect 497182 636392 497188 636404
rect 72476 636364 497188 636392
rect 72476 636352 72482 636364
rect 497182 636352 497188 636364
rect 497240 636352 497246 636404
rect 21358 636284 21364 636336
rect 21416 636324 21422 636336
rect 451918 636324 451924 636336
rect 21416 636296 451924 636324
rect 21416 636284 21422 636296
rect 451918 636284 451924 636296
rect 451976 636284 451982 636336
rect 94222 636216 94228 636268
rect 94280 636256 94286 636268
rect 531958 636256 531964 636268
rect 94280 636228 531964 636256
rect 94280 636216 94286 636228
rect 531958 636216 531964 636228
rect 532016 636216 532022 636268
rect 293862 635672 293868 635724
rect 293920 635712 293926 635724
rect 299474 635712 299480 635724
rect 293920 635684 299480 635712
rect 293920 635672 293926 635684
rect 299474 635672 299480 635684
rect 299532 635672 299538 635724
rect 282822 635604 282828 635656
rect 282880 635644 282886 635656
rect 364334 635644 364340 635656
rect 282880 635616 364340 635644
rect 282880 635604 282886 635616
rect 364334 635604 364340 635616
rect 364392 635604 364398 635656
rect 271506 635536 271512 635588
rect 271564 635576 271570 635588
rect 429194 635576 429200 635588
rect 271564 635548 429200 635576
rect 271564 635536 271570 635548
rect 429194 635536 429200 635548
rect 429252 635536 429258 635588
rect 260190 635468 260196 635520
rect 260248 635508 260254 635520
rect 494054 635508 494060 635520
rect 260248 635480 494060 635508
rect 260248 635468 260254 635480
rect 494054 635468 494060 635480
rect 494112 635468 494118 635520
rect 226242 635400 226248 635452
rect 226300 635440 226306 635452
rect 512822 635440 512828 635452
rect 226300 635412 512828 635440
rect 226300 635400 226306 635412
rect 512822 635400 512828 635412
rect 512880 635400 512886 635452
rect 214926 635332 214932 635384
rect 214984 635372 214990 635384
rect 512730 635372 512736 635384
rect 214984 635344 512736 635372
rect 214984 635332 214990 635344
rect 512730 635332 512736 635344
rect 512788 635332 512794 635384
rect 71314 635264 71320 635316
rect 71372 635304 71378 635316
rect 372706 635304 372712 635316
rect 71372 635276 372712 635304
rect 71372 635264 71378 635276
rect 372706 635264 372712 635276
rect 372764 635264 372770 635316
rect 203610 635196 203616 635248
rect 203668 635236 203674 635248
rect 514294 635236 514300 635248
rect 203668 635208 514300 635236
rect 203668 635196 203674 635208
rect 514294 635196 514300 635208
rect 514352 635196 514358 635248
rect 71222 635128 71228 635180
rect 71280 635168 71286 635180
rect 384022 635168 384028 635180
rect 71280 635140 384028 635168
rect 71280 635128 71286 635140
rect 384022 635128 384028 635140
rect 384080 635128 384086 635180
rect 199838 635060 199844 635112
rect 199896 635100 199902 635112
rect 525242 635100 525248 635112
rect 199896 635072 525248 635100
rect 199896 635060 199902 635072
rect 525242 635060 525248 635072
rect 525300 635060 525306 635112
rect 62758 634992 62764 635044
rect 62816 635032 62822 635044
rect 395338 635032 395344 635044
rect 62816 635004 395344 635032
rect 62816 634992 62822 635004
rect 395338 634992 395344 635004
rect 395396 634992 395402 635044
rect 71130 634924 71136 634976
rect 71188 634964 71194 634976
rect 406654 634964 406660 634976
rect 71188 634936 406660 634964
rect 71188 634924 71194 634936
rect 406654 634924 406660 634936
rect 406712 634924 406718 634976
rect 3510 634856 3516 634908
rect 3568 634896 3574 634908
rect 361574 634896 361580 634908
rect 3568 634868 361580 634896
rect 3568 634856 3574 634868
rect 361574 634856 361580 634868
rect 361632 634856 361638 634908
rect 113082 634788 113088 634840
rect 113140 634828 113146 634840
rect 514110 634828 514116 634840
rect 113140 634800 514116 634828
rect 113140 634788 113146 634800
rect 514110 634788 514116 634800
rect 514168 634788 514174 634840
rect 216674 634312 216680 634364
rect 216732 634352 216738 634364
rect 433426 634352 433432 634364
rect 216732 634324 433432 634352
rect 216732 634312 216738 634324
rect 433426 634312 433432 634324
rect 433484 634312 433490 634364
rect 139302 634244 139308 634296
rect 139360 634284 139366 634296
rect 365622 634284 365628 634296
rect 139360 634256 365628 634284
rect 139360 634244 139366 634256
rect 365622 634244 365628 634256
rect 365680 634244 365686 634296
rect 366542 634244 366548 634296
rect 366600 634284 366606 634296
rect 459554 634284 459560 634296
rect 366600 634256 459560 634284
rect 366600 634244 366606 634256
rect 459554 634244 459560 634256
rect 459612 634244 459618 634296
rect 177206 634176 177212 634228
rect 177264 634216 177270 634228
rect 525150 634216 525156 634228
rect 177264 634188 525156 634216
rect 177264 634176 177270 634188
rect 525150 634176 525156 634188
rect 525208 634176 525214 634228
rect 192294 634108 192300 634160
rect 192352 634148 192358 634160
rect 545758 634148 545764 634160
rect 192352 634120 545764 634148
rect 192352 634108 192358 634120
rect 545758 634108 545764 634120
rect 545816 634108 545822 634160
rect 165890 634040 165896 634092
rect 165948 634080 165954 634092
rect 525058 634080 525064 634092
rect 165948 634052 525064 634080
rect 165948 634040 165954 634052
rect 525058 634040 525064 634052
rect 525116 634040 525122 634092
rect 154482 633972 154488 634024
rect 154540 634012 154546 634024
rect 522298 634012 522304 634024
rect 154540 633984 522304 634012
rect 154540 633972 154546 633984
rect 522298 633972 522304 633984
rect 522356 633972 522362 634024
rect 131942 633904 131948 633956
rect 132000 633944 132006 633956
rect 518158 633944 518164 633956
rect 132000 633916 518164 633944
rect 132000 633904 132006 633916
rect 518158 633904 518164 633916
rect 518216 633904 518222 633956
rect 4062 633836 4068 633888
rect 4120 633876 4126 633888
rect 391934 633876 391940 633888
rect 4120 633848 391940 633876
rect 4120 633836 4126 633848
rect 391934 633836 391940 633848
rect 391992 633836 391998 633888
rect 3878 633768 3884 633820
rect 3936 633808 3942 633820
rect 425514 633808 425520 633820
rect 3936 633780 425520 633808
rect 3936 633768 3942 633780
rect 425514 633768 425520 633780
rect 425572 633768 425578 633820
rect 3786 633700 3792 633752
rect 3844 633740 3850 633752
rect 436830 633740 436836 633752
rect 3844 633712 436836 633740
rect 3844 633700 3850 633712
rect 436830 633700 436836 633712
rect 436888 633700 436894 633752
rect 4982 633632 4988 633684
rect 5040 633672 5046 633684
rect 448514 633672 448520 633684
rect 5040 633644 448520 633672
rect 5040 633632 5046 633644
rect 448514 633632 448520 633644
rect 448572 633632 448578 633684
rect 3418 633564 3424 633616
rect 3476 633604 3482 633616
rect 455690 633604 455696 633616
rect 3476 633576 455696 633604
rect 3476 633564 3482 633576
rect 455690 633564 455696 633576
rect 455748 633564 455754 633616
rect 505370 633564 505376 633616
rect 505428 633604 505434 633616
rect 511994 633604 512000 633616
rect 505428 633576 512000 633604
rect 505428 633564 505434 633576
rect 511994 633564 512000 633576
rect 512052 633564 512058 633616
rect 4890 633496 4896 633548
rect 4948 633536 4954 633548
rect 470870 633536 470876 633548
rect 4948 633508 470876 633536
rect 4948 633496 4954 633508
rect 470870 633496 470876 633508
rect 470928 633496 470934 633548
rect 501598 633496 501604 633548
rect 501656 633536 501662 633548
rect 511074 633536 511080 633548
rect 501656 633508 511080 633536
rect 501656 633496 501662 633508
rect 511074 633496 511080 633508
rect 511132 633496 511138 633548
rect 4798 633428 4804 633480
rect 4856 633468 4862 633480
rect 482094 633468 482100 633480
rect 4856 633440 482100 633468
rect 4856 633428 4862 633440
rect 482094 633428 482100 633440
rect 482152 633428 482158 633480
rect 493962 633428 493968 633480
rect 494020 633468 494026 633480
rect 512086 633468 512092 633480
rect 494020 633440 512092 633468
rect 494020 633428 494026 633440
rect 512086 633428 512092 633440
rect 512144 633428 512150 633480
rect 5258 632884 5264 632936
rect 5316 632924 5322 632936
rect 365162 632924 365168 632936
rect 5316 632896 365168 632924
rect 5316 632884 5322 632896
rect 365162 632884 365168 632896
rect 365220 632884 365226 632936
rect 158346 632816 158352 632868
rect 158404 632856 158410 632868
rect 511442 632856 511448 632868
rect 158404 632828 511448 632856
rect 158404 632816 158410 632828
rect 511442 632816 511448 632828
rect 511500 632816 511506 632868
rect 3694 632748 3700 632800
rect 3752 632788 3758 632800
rect 216674 632788 216680 632800
rect 3752 632760 216680 632788
rect 3752 632748 3758 632760
rect 216674 632748 216680 632760
rect 216732 632748 216738 632800
rect 222470 632748 222476 632800
rect 222528 632788 222534 632800
rect 579982 632788 579988 632800
rect 222528 632760 579988 632788
rect 222528 632748 222534 632760
rect 579982 632748 579988 632760
rect 580040 632748 580046 632800
rect 365622 632680 365628 632732
rect 365680 632720 365686 632732
rect 580442 632720 580448 632732
rect 365680 632692 580448 632720
rect 365680 632680 365686 632692
rect 580442 632680 580448 632692
rect 580500 632680 580506 632732
rect 218698 632612 218704 632664
rect 218756 632652 218762 632664
rect 580074 632652 580080 632664
rect 218756 632624 580080 632652
rect 218756 632612 218762 632624
rect 580074 632612 580080 632624
rect 580132 632612 580138 632664
rect 3326 632544 3332 632596
rect 3384 632584 3390 632596
rect 376846 632584 376852 632596
rect 3384 632556 376852 632584
rect 3384 632544 3390 632556
rect 376846 632544 376852 632556
rect 376904 632544 376910 632596
rect 207382 632476 207388 632528
rect 207440 632516 207446 632528
rect 580902 632516 580908 632528
rect 207440 632488 580908 632516
rect 207440 632476 207446 632488
rect 580902 632476 580908 632488
rect 580960 632476 580966 632528
rect 135714 632408 135720 632460
rect 135772 632448 135778 632460
rect 511350 632448 511356 632460
rect 135772 632420 511356 632448
rect 135772 632408 135778 632420
rect 511350 632408 511356 632420
rect 511408 632408 511414 632460
rect 3234 632340 3240 632392
rect 3292 632380 3298 632392
rect 380250 632380 380256 632392
rect 3292 632352 380256 632380
rect 3292 632340 3298 632352
rect 380250 632340 380256 632352
rect 380308 632340 380314 632392
rect 195882 632272 195888 632324
rect 195940 632312 195946 632324
rect 580718 632312 580724 632324
rect 195940 632284 580724 632312
rect 195940 632272 195946 632284
rect 580718 632272 580724 632284
rect 580776 632272 580782 632324
rect 3970 632204 3976 632256
rect 4028 632244 4034 632256
rect 399110 632244 399116 632256
rect 4028 632216 399116 632244
rect 4028 632204 4034 632216
rect 399110 632204 399116 632216
rect 399168 632204 399174 632256
rect 3602 632136 3608 632188
rect 3660 632176 3666 632188
rect 444696 632176 444702 632188
rect 3660 632148 444702 632176
rect 3660 632136 3666 632148
rect 444696 632136 444702 632148
rect 444754 632136 444760 632188
rect 127848 632068 127854 632120
rect 127906 632108 127912 632120
rect 580258 632108 580264 632120
rect 127906 632080 580264 632108
rect 127906 632068 127912 632080
rect 580258 632068 580264 632080
rect 580316 632068 580322 632120
rect 410058 631660 410064 631712
rect 410116 631700 410122 631712
rect 421006 631700 421012 631712
rect 410116 631672 421012 631700
rect 410116 631660 410122 631672
rect 421006 631660 421012 631672
rect 421064 631660 421070 631712
rect 408466 631604 425054 631632
rect 142798 631524 142804 631576
rect 142856 631564 142862 631576
rect 146938 631564 146944 631576
rect 142856 631536 146944 631564
rect 142856 631524 142862 631536
rect 146938 631524 146944 631536
rect 146996 631524 147002 631576
rect 135226 631468 150434 631496
rect 5166 630776 5172 630828
rect 5224 630816 5230 630828
rect 135226 630816 135254 631468
rect 142798 631428 142804 631440
rect 5224 630788 135254 630816
rect 142126 631400 142804 631428
rect 5224 630776 5230 630788
rect 5074 630708 5080 630760
rect 5132 630748 5138 630760
rect 5132 630720 136634 630748
rect 5132 630708 5138 630720
rect 136606 630408 136634 630720
rect 142126 630408 142154 631400
rect 142798 631388 142804 631400
rect 142856 631388 142862 631440
rect 143258 631388 143264 631440
rect 143316 631388 143322 631440
rect 146938 631388 146944 631440
rect 146996 631388 147002 631440
rect 136606 630380 142154 630408
rect 143276 630136 143304 631388
rect 146956 630816 146984 631388
rect 150406 630884 150434 631468
rect 169662 631388 169668 631440
rect 169720 631428 169726 631440
rect 169720 631400 171134 631428
rect 169720 631388 169726 631400
rect 171106 630884 171134 631400
rect 188522 631388 188528 631440
rect 188580 631428 188586 631440
rect 188580 631400 190454 631428
rect 188580 631388 188586 631400
rect 190426 630952 190454 631400
rect 211062 631388 211068 631440
rect 211120 631428 211126 631440
rect 211120 631400 219434 631428
rect 211120 631388 211126 631400
rect 219406 631020 219434 631400
rect 233786 631388 233792 631440
rect 233844 631428 233850 631440
rect 233844 631400 238754 631428
rect 233844 631388 233850 631400
rect 238726 631088 238754 631400
rect 408466 631088 408494 631604
rect 425026 631564 425054 631604
rect 410168 631536 416544 631564
rect 425026 631536 430574 631564
rect 410058 631388 410064 631440
rect 410116 631388 410122 631440
rect 238726 631060 408494 631088
rect 410076 631020 410104 631388
rect 219406 630992 410104 631020
rect 410168 630952 410196 631536
rect 190426 630924 410196 630952
rect 410260 631468 410656 631496
rect 410260 630884 410288 631468
rect 410518 631388 410524 631440
rect 410576 631388 410582 631440
rect 410536 631020 410564 631388
rect 410628 631360 410656 631468
rect 415366 631468 415900 631496
rect 415366 631428 415394 631468
rect 411226 631400 415394 631428
rect 411226 631360 411254 631400
rect 415486 631388 415492 631440
rect 415544 631388 415550 631440
rect 410628 631332 411254 631360
rect 415504 631088 415532 631388
rect 415872 631224 415900 631468
rect 416516 631360 416544 631536
rect 421006 631456 421012 631508
rect 421064 631496 421070 631508
rect 421064 631468 430160 631496
rect 421064 631456 421070 631468
rect 416590 631388 416596 631440
rect 416648 631428 416654 631440
rect 416648 631400 427814 631428
rect 416648 631388 416654 631400
rect 416516 631332 425054 631360
rect 415872 631196 418338 631224
rect 150406 630856 154574 630884
rect 171106 630856 410288 630884
rect 410444 630992 410564 631020
rect 415366 631060 415532 631088
rect 154546 630816 154574 630856
rect 410444 630816 410472 630992
rect 146956 630788 151814 630816
rect 154546 630788 410472 630816
rect 411226 630856 411484 630884
rect 151786 630680 151814 630788
rect 411226 630748 411254 630856
rect 411456 630816 411484 630856
rect 415366 630816 415394 631060
rect 418310 630952 418338 631196
rect 425026 631020 425054 631332
rect 427786 631292 427814 631400
rect 429286 631388 429292 631440
rect 429344 631388 429350 631440
rect 429304 631292 429332 631388
rect 427786 631264 429332 631292
rect 430132 631020 430160 631468
rect 430546 631088 430574 631536
rect 580166 631088 580172 631100
rect 430546 631060 580172 631088
rect 580166 631048 580172 631060
rect 580224 631048 580230 631100
rect 580810 631020 580816 631032
rect 425026 630992 427814 631020
rect 430132 630992 580816 631020
rect 418310 630924 425054 630952
rect 411456 630788 415394 630816
rect 153166 630720 411254 630748
rect 153166 630680 153194 630720
rect 151786 630652 153194 630680
rect 154546 630652 411254 630680
rect 154546 630612 154574 630652
rect 153166 630584 154574 630612
rect 153166 630136 153194 630584
rect 411226 630408 411254 630652
rect 425026 630612 425054 630924
rect 427786 630884 427814 630992
rect 580810 630980 580816 630992
rect 580868 630980 580874 631032
rect 580626 630952 580632 630964
rect 431926 630924 580632 630952
rect 427786 630856 429424 630884
rect 429396 630816 429424 630856
rect 431926 630816 431954 630924
rect 580626 630912 580632 630924
rect 580684 630912 580690 630964
rect 580534 630884 580540 630896
rect 429396 630788 431954 630816
rect 434686 630856 580540 630884
rect 434686 630748 434714 630856
rect 580534 630844 580540 630856
rect 580592 630844 580598 630896
rect 429396 630720 434714 630748
rect 429396 630680 429424 630720
rect 579982 630708 579988 630760
rect 580040 630748 580046 630760
rect 580166 630748 580172 630760
rect 580040 630720 580172 630748
rect 580040 630708 580046 630720
rect 580166 630708 580172 630720
rect 580224 630708 580230 630760
rect 580350 630680 580356 630692
rect 429166 630652 429424 630680
rect 430546 630652 580356 630680
rect 429166 630612 429194 630652
rect 425026 630584 429194 630612
rect 430546 630408 430574 630652
rect 580350 630640 580356 630652
rect 580408 630640 580414 630692
rect 411226 630380 430574 630408
rect 143276 630108 153194 630136
rect 3142 619556 3148 619608
rect 3200 619596 3206 619608
rect 68370 619596 68376 619608
rect 3200 619568 68376 619596
rect 3200 619556 3206 619568
rect 68370 619556 68376 619568
rect 68428 619556 68434 619608
rect 512822 618196 512828 618248
rect 512880 618236 512886 618248
rect 579982 618236 579988 618248
rect 512880 618208 579988 618236
rect 512880 618196 512886 618208
rect 579982 618196 579988 618208
rect 580040 618196 580046 618248
rect 2774 607044 2780 607096
rect 2832 607084 2838 607096
rect 5258 607084 5264 607096
rect 2832 607056 5264 607084
rect 2832 607044 2838 607056
rect 5258 607044 5264 607056
rect 5316 607044 5322 607096
rect 3142 580932 3148 580984
rect 3200 580972 3206 580984
rect 71314 580972 71320 580984
rect 3200 580944 71320 580972
rect 3200 580932 3206 580944
rect 71314 580932 71320 580944
rect 71372 580932 71378 580984
rect 512730 564340 512736 564392
rect 512788 564380 512794 564392
rect 580166 564380 580172 564392
rect 512788 564352 580172 564380
rect 512788 564340 512794 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3326 528504 3332 528556
rect 3384 528544 3390 528556
rect 71222 528544 71228 528556
rect 3384 528516 71228 528544
rect 3384 528504 3390 528516
rect 71222 528504 71228 528516
rect 71280 528504 71286 528556
rect 514294 511912 514300 511964
rect 514352 511952 514358 511964
rect 580166 511952 580172 511964
rect 514352 511924 580172 511952
rect 514352 511912 514358 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3326 501780 3332 501832
rect 3384 501820 3390 501832
rect 7558 501820 7564 501832
rect 3384 501792 7564 501820
rect 3384 501780 3390 501792
rect 7558 501780 7564 501792
rect 7616 501780 7622 501832
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 62758 476048 62764 476060
rect 3384 476020 62764 476048
rect 3384 476008 3390 476020
rect 62758 476008 62764 476020
rect 62816 476008 62822 476060
rect 525242 471928 525248 471980
rect 525300 471968 525306 471980
rect 579798 471968 579804 471980
rect 525300 471940 579804 471968
rect 525300 471928 525306 471940
rect 579798 471928 579804 471940
rect 579856 471928 579862 471980
rect 3326 463632 3332 463684
rect 3384 463672 3390 463684
rect 58618 463672 58624 463684
rect 3384 463644 58624 463672
rect 3384 463632 3390 463644
rect 58618 463632 58624 463644
rect 58676 463632 58682 463684
rect 545758 458124 545764 458176
rect 545816 458164 545822 458176
rect 580166 458164 580172 458176
rect 545816 458136 580172 458164
rect 545816 458124 545822 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 522390 431876 522396 431928
rect 522448 431916 522454 431928
rect 580166 431916 580172 431928
rect 522448 431888 580172 431916
rect 522448 431876 522454 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 71130 423620 71136 423632
rect 3384 423592 71136 423620
rect 3384 423580 3390 423592
rect 71130 423580 71136 423592
rect 71188 423580 71194 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 53098 411244 53104 411256
rect 3384 411216 53104 411244
rect 3384 411204 3390 411216
rect 53098 411204 53104 411216
rect 53156 411204 53162 411256
rect 516962 405628 516968 405680
rect 517020 405668 517026 405680
rect 580166 405668 580172 405680
rect 517020 405640 580172 405668
rect 517020 405628 517026 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 13078 398800 13084 398812
rect 3384 398772 13084 398800
rect 3384 398760 3390 398772
rect 13078 398760 13084 398772
rect 13136 398760 13142 398812
rect 521010 379448 521016 379500
rect 521068 379488 521074 379500
rect 579614 379488 579620 379500
rect 521068 379460 579620 379488
rect 521068 379448 521074 379460
rect 579614 379448 579620 379460
rect 579672 379448 579678 379500
rect 2774 372308 2780 372360
rect 2832 372348 2838 372360
rect 5166 372348 5172 372360
rect 2832 372320 5172 372348
rect 2832 372308 2838 372320
rect 5166 372308 5172 372320
rect 5224 372308 5230 372360
rect 525150 365644 525156 365696
rect 525208 365684 525214 365696
rect 580166 365684 580172 365696
rect 525208 365656 580172 365684
rect 525208 365644 525214 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 2958 346332 2964 346384
rect 3016 346372 3022 346384
rect 57238 346372 57244 346384
rect 3016 346344 57244 346372
rect 3016 346332 3022 346344
rect 57238 346332 57244 346344
rect 57296 346332 57302 346384
rect 520918 325592 520924 325644
rect 520976 325632 520982 325644
rect 580166 325632 580172 325644
rect 520976 325604 580172 325632
rect 520976 325592 520982 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 2774 319812 2780 319864
rect 2832 319852 2838 319864
rect 5074 319852 5080 319864
rect 2832 319824 5080 319852
rect 2832 319812 2838 319824
rect 5074 319812 5080 319824
rect 5132 319812 5138 319864
rect 525058 313216 525064 313268
rect 525116 313256 525122 313268
rect 579706 313256 579712 313268
rect 525116 313228 579712 313256
rect 525116 313216 525122 313228
rect 579706 313216 579712 313228
rect 579764 313216 579770 313268
rect 511442 299412 511448 299464
rect 511500 299452 511506 299464
rect 579798 299452 579804 299464
rect 511500 299424 579804 299452
rect 511500 299412 511506 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 518250 273164 518256 273216
rect 518308 273204 518314 273216
rect 580166 273204 580172 273216
rect 518308 273176 580172 273204
rect 518308 273164 518314 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 66898 267696 66904 267708
rect 3292 267668 66904 267696
rect 3292 267656 3298 267668
rect 66898 267656 66904 267668
rect 66956 267656 66962 267708
rect 522298 259360 522304 259412
rect 522356 259400 522362 259412
rect 580166 259400 580172 259412
rect 522356 259372 580172 259400
rect 522356 259360 522362 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 2774 254940 2780 254992
rect 2832 254980 2838 254992
rect 4982 254980 4988 254992
rect 2832 254952 4988 254980
rect 2832 254940 2838 254952
rect 4982 254940 4988 254952
rect 5040 254940 5046 254992
rect 516870 245556 516876 245608
rect 516928 245596 516934 245608
rect 580166 245596 580172 245608
rect 516928 245568 580172 245596
rect 516928 245556 516934 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 21358 215268 21364 215280
rect 3384 215240 21364 215268
rect 3384 215228 3390 215240
rect 21358 215228 21364 215240
rect 21416 215228 21422 215280
rect 511350 206932 511356 206984
rect 511408 206972 511414 206984
rect 580166 206972 580172 206984
rect 511408 206944 580172 206972
rect 511408 206932 511414 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 518158 179324 518164 179376
rect 518216 179364 518222 179376
rect 580166 179364 580172 179376
rect 518216 179336 580172 179364
rect 518216 179324 518222 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 514202 166948 514208 167000
rect 514260 166988 514266 167000
rect 580166 166988 580172 167000
rect 514260 166960 580172 166988
rect 514260 166948 514266 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 71038 164200 71044 164212
rect 3292 164172 71044 164200
rect 3292 164160 3298 164172
rect 71038 164160 71044 164172
rect 71096 164160 71102 164212
rect 2774 149880 2780 149932
rect 2832 149920 2838 149932
rect 4890 149920 4896 149932
rect 2832 149892 4896 149920
rect 2832 149880 2838 149892
rect 4890 149880 4896 149892
rect 4948 149880 4954 149932
rect 514110 126896 514116 126948
rect 514168 126936 514174 126948
rect 580166 126936 580172 126948
rect 514168 126908 580172 126936
rect 514168 126896 514174 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 516778 113092 516784 113144
rect 516836 113132 516842 113144
rect 579798 113132 579804 113144
rect 516836 113104 579804 113132
rect 516836 113092 516842 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 64138 111772 64144 111784
rect 3476 111744 64144 111772
rect 3476 111732 3482 111744
rect 64138 111732 64144 111744
rect 64196 111732 64202 111784
rect 515398 100648 515404 100700
rect 515456 100688 515462 100700
rect 580166 100688 580172 100700
rect 515456 100660 580172 100688
rect 515456 100648 515462 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 511258 86912 511264 86964
rect 511316 86952 511322 86964
rect 580166 86952 580172 86964
rect 511316 86924 580172 86952
rect 511316 86912 511322 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 531958 73108 531964 73160
rect 532016 73148 532022 73160
rect 580166 73148 580172 73160
rect 532016 73120 580172 73148
rect 532016 73108 532022 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 89714 71884 89720 71936
rect 89772 71924 89778 71936
rect 90772 71924 90778 71936
rect 89772 71896 90778 71924
rect 89772 71884 89778 71896
rect 90772 71884 90778 71896
rect 90830 71884 90836 71936
rect 110414 71884 110420 71936
rect 110472 71924 110478 71936
rect 111472 71924 111478 71936
rect 110472 71896 111478 71924
rect 110472 71884 110478 71896
rect 111472 71884 111478 71896
rect 111530 71884 111536 71936
rect 114554 71884 114560 71936
rect 114612 71924 114618 71936
rect 115612 71924 115618 71936
rect 114612 71896 115618 71924
rect 114612 71884 114618 71896
rect 115612 71884 115618 71896
rect 115670 71884 115676 71936
rect 122834 71884 122840 71936
rect 122892 71924 122898 71936
rect 123892 71924 123898 71936
rect 122892 71896 123898 71924
rect 122892 71884 122898 71896
rect 123892 71884 123898 71896
rect 123950 71884 123956 71936
rect 131114 71884 131120 71936
rect 131172 71924 131178 71936
rect 132172 71924 132178 71936
rect 131172 71896 132178 71924
rect 131172 71884 131178 71896
rect 132172 71884 132178 71896
rect 132230 71884 132236 71936
rect 135254 71884 135260 71936
rect 135312 71924 135318 71936
rect 136312 71924 136318 71936
rect 135312 71896 136318 71924
rect 135312 71884 135318 71896
rect 136312 71884 136318 71896
rect 136370 71884 136376 71936
rect 147674 71884 147680 71936
rect 147732 71924 147738 71936
rect 148732 71924 148738 71936
rect 147732 71896 148738 71924
rect 147732 71884 147738 71896
rect 148732 71884 148738 71896
rect 148790 71884 148796 71936
rect 160094 71884 160100 71936
rect 160152 71924 160158 71936
rect 161152 71924 161158 71936
rect 160152 71896 161158 71924
rect 160152 71884 160158 71896
rect 161152 71884 161158 71896
rect 161210 71884 161216 71936
rect 176654 71884 176660 71936
rect 176712 71924 176718 71936
rect 177712 71924 177718 71936
rect 176712 71896 177718 71924
rect 176712 71884 176718 71896
rect 177712 71884 177718 71896
rect 177770 71884 177776 71936
rect 197446 71884 197452 71936
rect 197504 71924 197510 71936
rect 198412 71924 198418 71936
rect 197504 71896 198418 71924
rect 197504 71884 197510 71896
rect 198412 71884 198418 71896
rect 198470 71884 198476 71936
rect 201494 71884 201500 71936
rect 201552 71924 201558 71936
rect 202552 71924 202558 71936
rect 201552 71896 202558 71924
rect 201552 71884 201558 71896
rect 202552 71884 202558 71896
rect 202610 71884 202616 71936
rect 213914 71884 213920 71936
rect 213972 71924 213978 71936
rect 214972 71924 214978 71936
rect 213972 71896 214978 71924
rect 213972 71884 213978 71896
rect 214972 71884 214978 71896
rect 215030 71884 215036 71936
rect 296806 71884 296812 71936
rect 296864 71924 296870 71936
rect 297772 71924 297778 71936
rect 296864 71896 297778 71924
rect 296864 71884 296870 71896
rect 297772 71884 297778 71896
rect 297830 71884 297836 71936
rect 309134 71884 309140 71936
rect 309192 71924 309198 71936
rect 310192 71924 310198 71936
rect 309192 71896 310198 71924
rect 309192 71884 309198 71896
rect 310192 71884 310198 71896
rect 310250 71884 310256 71936
rect 346486 71884 346492 71936
rect 346544 71924 346550 71936
rect 347452 71924 347458 71936
rect 346544 71896 347458 71924
rect 346544 71884 346550 71896
rect 347452 71884 347458 71896
rect 347510 71884 347516 71936
rect 367094 71884 367100 71936
rect 367152 71924 367158 71936
rect 368152 71924 368158 71936
rect 367152 71896 368158 71924
rect 367152 71884 367158 71896
rect 368152 71884 368158 71896
rect 368210 71884 368216 71936
rect 412634 71884 412640 71936
rect 412692 71924 412698 71936
rect 413692 71924 413698 71936
rect 412692 71896 413698 71924
rect 412692 71884 412698 71896
rect 413692 71884 413698 71896
rect 413750 71884 413756 71936
rect 441614 71884 441620 71936
rect 441672 71924 441678 71936
rect 442672 71924 442678 71936
rect 441672 71896 442678 71924
rect 441672 71884 441678 71896
rect 442672 71884 442678 71896
rect 442730 71884 442736 71936
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 68278 71720 68284 71732
rect 3476 71692 68284 71720
rect 3476 71680 3482 71692
rect 68278 71680 68284 71692
rect 68336 71680 68342 71732
rect 233326 70320 233332 70372
rect 233384 70360 233390 70372
rect 251358 70360 251364 70372
rect 233384 70332 251364 70360
rect 233384 70320 233390 70332
rect 251358 70320 251364 70332
rect 251416 70320 251422 70372
rect 246298 70252 246304 70304
rect 246356 70292 246362 70304
rect 252186 70292 252192 70304
rect 246356 70264 252192 70292
rect 246356 70252 246362 70264
rect 252186 70252 252192 70264
rect 252244 70252 252250 70304
rect 77294 70184 77300 70236
rect 77352 70224 77358 70236
rect 142890 70224 142896 70236
rect 77352 70196 142896 70224
rect 77352 70184 77358 70196
rect 142890 70184 142896 70196
rect 142948 70184 142954 70236
rect 238018 70184 238024 70236
rect 238076 70224 238082 70236
rect 241514 70224 241520 70236
rect 238076 70196 241520 70224
rect 238076 70184 238082 70196
rect 241514 70184 241520 70196
rect 241572 70184 241578 70236
rect 247678 70184 247684 70236
rect 247736 70224 247742 70236
rect 254670 70224 254676 70236
rect 247736 70196 254676 70224
rect 247736 70184 247742 70196
rect 254670 70184 254676 70196
rect 254728 70184 254734 70236
rect 260834 70184 260840 70236
rect 260892 70224 260898 70236
rect 271230 70224 271236 70236
rect 260892 70196 271236 70224
rect 260892 70184 260898 70196
rect 271230 70184 271236 70196
rect 271288 70184 271294 70236
rect 494698 70224 494704 70236
rect 489886 70196 494704 70224
rect 50338 70116 50344 70168
rect 50396 70156 50402 70168
rect 118050 70156 118056 70168
rect 50396 70128 118056 70156
rect 50396 70116 50402 70128
rect 118050 70116 118056 70128
rect 118108 70116 118114 70168
rect 217318 70116 217324 70168
rect 217376 70156 217382 70168
rect 229094 70156 229100 70168
rect 217376 70128 229100 70156
rect 217376 70116 217382 70128
rect 229094 70116 229100 70128
rect 229152 70116 229158 70168
rect 256694 70116 256700 70168
rect 256752 70156 256758 70168
rect 267918 70156 267924 70168
rect 256752 70128 267924 70156
rect 256752 70116 256758 70128
rect 267918 70116 267924 70128
rect 267976 70116 267982 70168
rect 483290 70116 483296 70168
rect 483348 70156 483354 70168
rect 489886 70156 489914 70196
rect 494698 70184 494704 70196
rect 494756 70184 494762 70236
rect 494882 70184 494888 70236
rect 494940 70224 494946 70236
rect 549898 70224 549904 70236
rect 494940 70196 549904 70224
rect 494940 70184 494946 70196
rect 549898 70184 549904 70196
rect 549956 70184 549962 70236
rect 483348 70128 489914 70156
rect 483348 70116 483354 70128
rect 493226 70116 493232 70168
rect 493284 70156 493290 70168
rect 548518 70156 548524 70168
rect 493284 70128 548524 70156
rect 493284 70116 493290 70128
rect 548518 70116 548524 70128
rect 548576 70116 548582 70168
rect 70394 70048 70400 70100
rect 70452 70088 70458 70100
rect 138014 70088 138020 70100
rect 70452 70060 138020 70088
rect 70452 70048 70458 70060
rect 138014 70048 138020 70060
rect 138072 70048 138078 70100
rect 198734 70048 198740 70100
rect 198792 70088 198798 70100
rect 227346 70088 227352 70100
rect 198792 70060 227352 70088
rect 198792 70048 198798 70060
rect 227346 70048 227352 70060
rect 227404 70048 227410 70100
rect 254026 70048 254032 70100
rect 254084 70088 254090 70100
rect 266354 70088 266360 70100
rect 254084 70060 266360 70088
rect 254084 70048 254090 70060
rect 266354 70048 266360 70060
rect 266412 70048 266418 70100
rect 359090 70048 359096 70100
rect 359148 70088 359154 70100
rect 377398 70088 377404 70100
rect 359148 70060 377404 70088
rect 359148 70048 359154 70060
rect 377398 70048 377404 70060
rect 377456 70048 377462 70100
rect 416222 70048 416228 70100
rect 416280 70088 416286 70100
rect 450538 70088 450544 70100
rect 416280 70060 450544 70088
rect 416280 70048 416286 70060
rect 450538 70048 450544 70060
rect 450596 70048 450602 70100
rect 488258 70048 488264 70100
rect 488316 70088 488322 70100
rect 547138 70088 547144 70100
rect 488316 70060 489914 70088
rect 488316 70048 488322 70060
rect 39298 69980 39304 70032
rect 39356 70020 39362 70032
rect 113174 70020 113180 70032
rect 39356 69992 113180 70020
rect 39356 69980 39362 69992
rect 113174 69980 113180 69992
rect 113232 69980 113238 70032
rect 174538 69980 174544 70032
rect 174596 70020 174602 70032
rect 200114 70020 200120 70032
rect 174596 69992 200120 70020
rect 174596 69980 174602 69992
rect 200114 69980 200120 69992
rect 200172 69980 200178 70032
rect 221458 69980 221464 70032
rect 221516 70020 221522 70032
rect 233970 70020 233976 70032
rect 221516 69992 233976 70020
rect 221516 69980 221522 69992
rect 233970 69980 233976 69992
rect 234028 69980 234034 70032
rect 248414 69980 248420 70032
rect 248472 70020 248478 70032
rect 262214 70020 262220 70032
rect 248472 69992 262220 70020
rect 248472 69980 248478 69992
rect 262214 69980 262220 69992
rect 262272 69980 262278 70032
rect 263594 69980 263600 70032
rect 263652 70020 263658 70032
rect 272886 70020 272892 70032
rect 263652 69992 272892 70020
rect 263652 69980 263658 69992
rect 272886 69980 272892 69992
rect 272944 69980 272950 70032
rect 273254 69980 273260 70032
rect 273312 70020 273318 70032
rect 279510 70020 279516 70032
rect 273312 69992 279516 70020
rect 273312 69980 273318 69992
rect 279510 69980 279516 69992
rect 279568 69980 279574 70032
rect 361574 69980 361580 70032
rect 361632 70020 361638 70032
rect 382918 70020 382924 70032
rect 361632 69992 382924 70020
rect 361632 69980 361638 69992
rect 382918 69980 382924 69992
rect 382976 69980 382982 70032
rect 408770 69980 408776 70032
rect 408828 70020 408834 70032
rect 443638 70020 443644 70032
rect 408828 69992 443644 70020
rect 408828 69980 408834 69992
rect 443638 69980 443644 69992
rect 443696 69980 443702 70032
rect 465902 69980 465908 70032
rect 465960 70020 465966 70032
rect 478138 70020 478144 70032
rect 465960 69992 478144 70020
rect 465960 69980 465966 69992
rect 478138 69980 478144 69992
rect 478196 69980 478202 70032
rect 489886 70020 489914 70060
rect 493244 70060 547144 70088
rect 493244 70020 493272 70060
rect 547138 70048 547144 70060
rect 547196 70048 547202 70100
rect 489886 69992 493272 70020
rect 494698 69980 494704 70032
rect 494756 70020 494762 70032
rect 545758 70020 545764 70032
rect 494756 69992 545764 70020
rect 494756 69980 494762 69992
rect 545758 69980 545764 69992
rect 545816 69980 545822 70032
rect 28258 69912 28264 69964
rect 28316 69952 28322 69964
rect 102318 69952 102324 69964
rect 28316 69924 102324 69952
rect 28316 69912 28322 69924
rect 102318 69912 102324 69924
rect 102376 69912 102382 69964
rect 135898 69912 135904 69964
rect 135956 69952 135962 69964
rect 145374 69952 145380 69964
rect 135956 69924 145380 69952
rect 135956 69912 135962 69924
rect 145374 69912 145380 69924
rect 145432 69912 145438 69964
rect 197354 69912 197360 69964
rect 197412 69952 197418 69964
rect 226518 69952 226524 69964
rect 197412 69924 226524 69952
rect 197412 69912 197418 69924
rect 226518 69912 226524 69924
rect 226576 69912 226582 69964
rect 228358 69912 228364 69964
rect 228416 69952 228422 69964
rect 246390 69952 246396 69964
rect 228416 69924 246396 69952
rect 228416 69912 228422 69924
rect 246390 69912 246396 69924
rect 246448 69912 246454 69964
rect 247034 69912 247040 69964
rect 247092 69952 247098 69964
rect 261294 69952 261300 69964
rect 247092 69924 261300 69952
rect 247092 69912 247098 69924
rect 261294 69912 261300 69924
rect 261352 69912 261358 69964
rect 266354 69912 266360 69964
rect 266412 69952 266418 69964
rect 274634 69952 274640 69964
rect 266412 69924 274640 69952
rect 266412 69912 266418 69924
rect 274634 69912 274640 69924
rect 274692 69912 274698 69964
rect 320174 69912 320180 69964
rect 320232 69952 320238 69964
rect 327718 69952 327724 69964
rect 320232 69924 327724 69952
rect 320232 69912 320238 69924
rect 327718 69912 327724 69924
rect 327776 69912 327782 69964
rect 373994 69912 374000 69964
rect 374052 69952 374058 69964
rect 398098 69952 398104 69964
rect 374052 69924 398104 69952
rect 374052 69912 374058 69924
rect 398098 69912 398104 69924
rect 398156 69912 398162 69964
rect 421190 69912 421196 69964
rect 421248 69952 421254 69964
rect 474734 69952 474740 69964
rect 421248 69924 474740 69952
rect 421248 69912 421254 69924
rect 474734 69912 474740 69924
rect 474792 69912 474798 69964
rect 478322 69912 478328 69964
rect 478380 69952 478386 69964
rect 542998 69952 543004 69964
rect 478380 69924 543004 69952
rect 478380 69912 478386 69924
rect 542998 69912 543004 69924
rect 543056 69912 543062 69964
rect 32398 69844 32404 69896
rect 32456 69884 32462 69896
rect 108114 69884 108120 69896
rect 32456 69856 108120 69884
rect 32456 69844 32462 69856
rect 108114 69844 108120 69856
rect 108172 69844 108178 69896
rect 140038 69844 140044 69896
rect 140096 69884 140102 69896
rect 150434 69884 150440 69896
rect 140096 69856 150440 69884
rect 140096 69844 140102 69856
rect 150434 69844 150440 69856
rect 150492 69844 150498 69896
rect 167638 69844 167644 69896
rect 167696 69884 167702 69896
rect 172514 69884 172520 69896
rect 167696 69856 172520 69884
rect 167696 69844 167702 69856
rect 172514 69844 172520 69856
rect 172572 69844 172578 69896
rect 191834 69844 191840 69896
rect 191892 69884 191898 69896
rect 222378 69884 222384 69896
rect 191892 69856 222384 69884
rect 191892 69844 191898 69856
rect 222378 69844 222384 69856
rect 222436 69844 222442 69896
rect 225598 69844 225604 69896
rect 225656 69884 225662 69896
rect 229830 69884 229836 69896
rect 225656 69856 229836 69884
rect 225656 69844 225662 69856
rect 229830 69844 229836 69856
rect 229888 69844 229894 69896
rect 235258 69844 235264 69896
rect 235316 69884 235322 69896
rect 239766 69884 239772 69896
rect 235316 69856 239772 69884
rect 235316 69844 235322 69856
rect 239766 69844 239772 69856
rect 239824 69844 239830 69896
rect 251266 69844 251272 69896
rect 251324 69884 251330 69896
rect 263778 69884 263784 69896
rect 251324 69856 263784 69884
rect 251324 69844 251330 69856
rect 263778 69844 263784 69856
rect 263836 69844 263842 69896
rect 264974 69844 264980 69896
rect 265032 69884 265038 69896
rect 273714 69884 273720 69896
rect 265032 69856 273720 69884
rect 265032 69844 265038 69856
rect 273714 69844 273720 69856
rect 273772 69844 273778 69896
rect 273898 69844 273904 69896
rect 273956 69884 273962 69896
rect 278774 69884 278780 69896
rect 273956 69856 278780 69884
rect 273956 69844 273962 69856
rect 278774 69844 278780 69856
rect 278832 69844 278838 69896
rect 306098 69844 306104 69896
rect 306156 69884 306162 69896
rect 307018 69884 307024 69896
rect 306156 69856 307024 69884
rect 306156 69844 306162 69856
rect 307018 69844 307024 69856
rect 307076 69844 307082 69896
rect 334250 69844 334256 69896
rect 334308 69884 334314 69896
rect 335998 69884 336004 69896
rect 334308 69856 336004 69884
rect 334308 69844 334314 69856
rect 335998 69844 336004 69856
rect 336056 69844 336062 69896
rect 350810 69844 350816 69896
rect 350868 69884 350874 69896
rect 355318 69884 355324 69896
rect 350868 69856 355324 69884
rect 350868 69844 350874 69856
rect 355318 69844 355324 69856
rect 355376 69844 355382 69896
rect 374638 69884 374644 69896
rect 364306 69856 374644 69884
rect 25498 69776 25504 69828
rect 25556 69816 25562 69828
rect 101490 69816 101496 69828
rect 25556 69788 101496 69816
rect 25556 69776 25562 69788
rect 101490 69776 101496 69788
rect 101548 69776 101554 69828
rect 144178 69776 144184 69828
rect 144236 69816 144242 69828
rect 155310 69816 155316 69828
rect 144236 69788 155316 69816
rect 144236 69776 144242 69788
rect 155310 69776 155316 69788
rect 155368 69776 155374 69828
rect 156598 69776 156604 69828
rect 156656 69816 156662 69828
rect 167730 69816 167736 69828
rect 156656 69788 167736 69816
rect 156656 69776 156662 69788
rect 167730 69776 167736 69788
rect 167788 69776 167794 69828
rect 170398 69776 170404 69828
rect 170456 69816 170462 69828
rect 204990 69816 204996 69828
rect 170456 69788 204996 69816
rect 170456 69776 170462 69788
rect 204990 69776 204996 69788
rect 205048 69776 205054 69828
rect 205634 69776 205640 69828
rect 205692 69816 205698 69828
rect 232314 69816 232320 69828
rect 205692 69788 232320 69816
rect 205692 69776 205698 69788
rect 232314 69776 232320 69788
rect 232372 69776 232378 69828
rect 235994 69776 236000 69828
rect 236052 69816 236058 69828
rect 253934 69816 253940 69828
rect 236052 69788 253940 69816
rect 236052 69776 236058 69788
rect 253934 69776 253940 69788
rect 253992 69776 253998 69828
rect 255314 69776 255320 69828
rect 255372 69816 255378 69828
rect 267090 69816 267096 69828
rect 255372 69788 267096 69816
rect 255372 69776 255378 69788
rect 267090 69776 267096 69788
rect 267148 69776 267154 69828
rect 285674 69776 285680 69828
rect 285732 69816 285738 69828
rect 288618 69816 288624 69828
rect 285732 69788 288624 69816
rect 285732 69776 285738 69788
rect 288618 69776 288624 69788
rect 288676 69776 288682 69828
rect 354122 69776 354128 69828
rect 354180 69816 354186 69828
rect 364306 69816 364334 69856
rect 374638 69844 374644 69856
rect 374696 69844 374702 69896
rect 376478 69844 376484 69896
rect 376536 69884 376542 69896
rect 400858 69884 400864 69896
rect 376536 69856 400864 69884
rect 376536 69844 376542 69856
rect 400858 69844 400864 69856
rect 400916 69844 400922 69896
rect 411254 69844 411260 69896
rect 411312 69884 411318 69896
rect 446398 69884 446404 69896
rect 411312 69856 446404 69884
rect 411312 69844 411318 69856
rect 446398 69844 446404 69856
rect 446456 69844 446462 69896
rect 453482 69844 453488 69896
rect 453540 69884 453546 69896
rect 521654 69884 521660 69896
rect 453540 69856 521660 69884
rect 453540 69844 453546 69856
rect 521654 69844 521660 69856
rect 521712 69844 521718 69896
rect 354180 69788 364334 69816
rect 354180 69776 354186 69788
rect 369026 69776 369032 69828
rect 369084 69816 369090 69828
rect 393958 69816 393964 69828
rect 369084 69788 393964 69816
rect 369084 69776 369090 69788
rect 393958 69776 393964 69788
rect 394016 69776 394022 69828
rect 403802 69776 403808 69828
rect 403860 69816 403866 69828
rect 440878 69816 440884 69828
rect 403860 69788 440884 69816
rect 403860 69776 403866 69788
rect 440878 69776 440884 69788
rect 440936 69776 440942 69828
rect 445754 69776 445760 69828
rect 445812 69816 445818 69828
rect 453298 69816 453304 69828
rect 445812 69788 453304 69816
rect 445812 69776 445818 69788
rect 453298 69776 453304 69788
rect 453356 69776 453362 69828
rect 458450 69776 458456 69828
rect 458508 69816 458514 69828
rect 528554 69816 528560 69828
rect 458508 69788 528560 69816
rect 458508 69776 458514 69788
rect 528554 69776 528560 69788
rect 528612 69776 528618 69828
rect 14458 69708 14464 69760
rect 14516 69748 14522 69760
rect 95694 69748 95700 69760
rect 14516 69720 95700 69748
rect 14516 69708 14522 69720
rect 95694 69708 95700 69720
rect 95752 69708 95758 69760
rect 124214 69708 124220 69760
rect 124272 69748 124278 69760
rect 175274 69748 175280 69760
rect 124272 69720 175280 69748
rect 124272 69708 124278 69720
rect 175274 69708 175280 69720
rect 175332 69708 175338 69760
rect 184934 69708 184940 69760
rect 184992 69748 184998 69760
rect 217410 69748 217416 69760
rect 184992 69720 217416 69748
rect 184992 69708 184998 69720
rect 217410 69708 217416 69720
rect 217468 69708 217474 69760
rect 229094 69708 229100 69760
rect 229152 69748 229158 69760
rect 248874 69748 248880 69760
rect 229152 69720 248880 69748
rect 229152 69708 229158 69720
rect 248874 69708 248880 69720
rect 248932 69708 248938 69760
rect 251174 69708 251180 69760
rect 251232 69748 251238 69760
rect 264606 69748 264612 69760
rect 251232 69720 264612 69748
rect 251232 69708 251238 69720
rect 264606 69708 264612 69720
rect 264664 69708 264670 69760
rect 335906 69708 335912 69760
rect 335964 69748 335970 69760
rect 345658 69748 345664 69760
rect 335964 69720 345664 69748
rect 335964 69708 335970 69720
rect 345658 69708 345664 69720
rect 345716 69708 345722 69760
rect 349154 69708 349160 69760
rect 349212 69748 349218 69760
rect 362218 69748 362224 69760
rect 349212 69720 362224 69748
rect 349212 69708 349218 69720
rect 362218 69708 362224 69720
rect 362276 69708 362282 69760
rect 385034 69748 385040 69760
rect 362328 69720 385040 69748
rect 10318 69640 10324 69692
rect 10376 69680 10382 69692
rect 91554 69680 91560 69692
rect 10376 69652 91560 69680
rect 10376 69640 10382 69652
rect 91554 69640 91560 69652
rect 91612 69640 91618 69692
rect 106274 69640 106280 69692
rect 106332 69680 106338 69692
rect 162854 69680 162860 69692
rect 106332 69652 162860 69680
rect 106332 69640 106338 69652
rect 162854 69640 162860 69652
rect 162912 69640 162918 69692
rect 169754 69640 169760 69692
rect 169812 69680 169818 69692
rect 207474 69680 207480 69692
rect 169812 69652 207480 69680
rect 169812 69640 169818 69652
rect 207474 69640 207480 69652
rect 207532 69640 207538 69692
rect 219434 69640 219440 69692
rect 219492 69680 219498 69692
rect 242250 69680 242256 69692
rect 219492 69652 242256 69680
rect 219492 69640 219498 69652
rect 242250 69640 242256 69652
rect 242308 69640 242314 69692
rect 242894 69640 242900 69692
rect 242952 69680 242958 69692
rect 258810 69680 258816 69692
rect 242952 69652 258816 69680
rect 242952 69640 242958 69652
rect 258810 69640 258816 69652
rect 258868 69640 258874 69692
rect 259454 69640 259460 69692
rect 259512 69680 259518 69692
rect 270494 69680 270500 69692
rect 259512 69652 270500 69680
rect 259512 69640 259518 69652
rect 270494 69640 270500 69652
rect 270552 69640 270558 69692
rect 274634 69640 274640 69692
rect 274692 69680 274698 69692
rect 280338 69680 280344 69692
rect 274692 69652 280344 69680
rect 274692 69640 274698 69652
rect 280338 69640 280344 69652
rect 280396 69640 280402 69692
rect 311894 69640 311900 69692
rect 311952 69680 311958 69692
rect 318794 69680 318800 69692
rect 311952 69652 318800 69680
rect 311952 69640 311958 69652
rect 318794 69640 318800 69652
rect 318852 69640 318858 69692
rect 325970 69640 325976 69692
rect 326028 69680 326034 69692
rect 336090 69680 336096 69692
rect 326028 69652 336096 69680
rect 326028 69640 326034 69652
rect 336090 69640 336096 69652
rect 336148 69640 336154 69692
rect 344186 69640 344192 69692
rect 344244 69680 344250 69692
rect 358078 69680 358084 69692
rect 344244 69652 358084 69680
rect 344244 69640 344250 69652
rect 358078 69640 358084 69652
rect 358136 69640 358142 69692
rect 358262 69640 358268 69692
rect 358320 69680 358326 69692
rect 362328 69680 362356 69720
rect 385034 69708 385040 69720
rect 385092 69708 385098 69760
rect 398834 69708 398840 69760
rect 398892 69748 398898 69760
rect 436738 69748 436744 69760
rect 398892 69720 436744 69748
rect 398892 69708 398898 69720
rect 436738 69708 436744 69720
rect 436796 69708 436802 69760
rect 468386 69708 468392 69760
rect 468444 69748 468450 69760
rect 540238 69748 540244 69760
rect 468444 69720 540244 69748
rect 468444 69708 468450 69720
rect 540238 69708 540244 69720
rect 540296 69708 540302 69760
rect 358320 69652 362356 69680
rect 358320 69640 358326 69652
rect 364058 69640 364064 69692
rect 364116 69680 364122 69692
rect 391198 69680 391204 69692
rect 364116 69652 391204 69680
rect 364116 69640 364122 69652
rect 391198 69640 391204 69652
rect 391256 69640 391262 69692
rect 393866 69640 393872 69692
rect 393924 69680 393930 69692
rect 435358 69680 435364 69692
rect 393924 69652 435364 69680
rect 393924 69640 393930 69652
rect 435358 69640 435364 69652
rect 435416 69640 435422 69692
rect 448514 69640 448520 69692
rect 448572 69680 448578 69692
rect 456058 69680 456064 69692
rect 448572 69652 456064 69680
rect 448572 69640 448578 69652
rect 456058 69640 456064 69652
rect 456116 69640 456122 69692
rect 463418 69640 463424 69692
rect 463476 69680 463482 69692
rect 535454 69680 535460 69692
rect 463476 69652 535460 69680
rect 463476 69640 463482 69652
rect 535454 69640 535460 69652
rect 535512 69640 535518 69692
rect 233878 69504 233884 69556
rect 233936 69544 233942 69556
rect 238938 69544 238944 69556
rect 233936 69516 238944 69544
rect 233936 69504 233942 69516
rect 238938 69504 238944 69516
rect 238996 69504 239002 69556
rect 242250 69504 242256 69556
rect 242308 69544 242314 69556
rect 249794 69544 249800 69556
rect 242308 69516 249800 69544
rect 242308 69504 242314 69516
rect 249794 69504 249800 69516
rect 249852 69504 249858 69556
rect 270494 69504 270500 69556
rect 270552 69544 270558 69556
rect 277854 69544 277860 69556
rect 270552 69516 277860 69544
rect 270552 69504 270558 69516
rect 277854 69504 277860 69516
rect 277912 69504 277918 69556
rect 267734 69300 267740 69352
rect 267792 69340 267798 69352
rect 276198 69340 276204 69352
rect 267792 69312 276204 69340
rect 267792 69300 267798 69312
rect 276198 69300 276204 69312
rect 276256 69300 276262 69352
rect 261478 69232 261484 69284
rect 261536 69272 261542 69284
rect 268746 69272 268752 69284
rect 261536 69244 268752 69272
rect 261536 69232 261542 69244
rect 268746 69232 268752 69244
rect 268804 69232 268810 69284
rect 277394 69232 277400 69284
rect 277452 69272 277458 69284
rect 282914 69272 282920 69284
rect 277452 69244 282920 69272
rect 277452 69232 277458 69244
rect 282914 69232 282920 69244
rect 282972 69232 282978 69284
rect 284294 69232 284300 69284
rect 284352 69272 284358 69284
rect 287790 69272 287796 69284
rect 284352 69244 287796 69272
rect 284352 69232 284358 69244
rect 287790 69232 287796 69244
rect 287848 69232 287854 69284
rect 300854 69232 300860 69284
rect 300912 69272 300918 69284
rect 303614 69272 303620 69284
rect 300912 69244 303620 69272
rect 300912 69232 300918 69244
rect 303614 69232 303620 69244
rect 303672 69232 303678 69284
rect 267826 69164 267832 69216
rect 267884 69204 267890 69216
rect 275370 69204 275376 69216
rect 267884 69176 275376 69204
rect 267884 69164 267890 69176
rect 275370 69164 275376 69176
rect 275428 69164 275434 69216
rect 280154 69164 280160 69216
rect 280212 69204 280218 69216
rect 284478 69204 284484 69216
rect 280212 69176 284484 69204
rect 280212 69164 280218 69176
rect 284478 69164 284484 69176
rect 284536 69164 284542 69216
rect 164878 69096 164884 69148
rect 164936 69136 164942 69148
rect 170214 69136 170220 69148
rect 164936 69108 170220 69136
rect 164936 69096 164942 69108
rect 170214 69096 170220 69108
rect 170272 69096 170278 69148
rect 239398 69096 239404 69148
rect 239456 69136 239462 69148
rect 247218 69136 247224 69148
rect 239456 69108 247224 69136
rect 239456 69096 239462 69108
rect 247218 69096 247224 69108
rect 247276 69096 247282 69148
rect 269114 69096 269120 69148
rect 269172 69136 269178 69148
rect 277026 69136 277032 69148
rect 269172 69108 277032 69136
rect 269172 69096 269178 69108
rect 277026 69096 277032 69108
rect 277084 69096 277090 69148
rect 278038 69096 278044 69148
rect 278096 69136 278102 69148
rect 281166 69136 281172 69148
rect 278096 69108 281172 69136
rect 278096 69096 278102 69108
rect 281166 69096 281172 69108
rect 281224 69096 281230 69148
rect 281534 69096 281540 69148
rect 281592 69136 281598 69148
rect 285306 69136 285312 69148
rect 281592 69108 285312 69136
rect 281592 69096 281598 69108
rect 285306 69096 285312 69108
rect 285364 69096 285370 69148
rect 287054 69096 287060 69148
rect 287112 69136 287118 69148
rect 289446 69136 289452 69148
rect 287112 69108 289452 69136
rect 287112 69096 287118 69108
rect 289446 69096 289452 69108
rect 289504 69096 289510 69148
rect 299474 69096 299480 69148
rect 299532 69136 299538 69148
rect 300854 69136 300860 69148
rect 299532 69108 300860 69136
rect 299532 69096 299538 69108
rect 300854 69096 300860 69108
rect 300912 69096 300918 69148
rect 308582 69096 308588 69148
rect 308640 69136 308646 69148
rect 311158 69136 311164 69148
rect 308640 69108 311164 69136
rect 308640 69096 308646 69108
rect 311158 69096 311164 69108
rect 311216 69096 311222 69148
rect 317690 69096 317696 69148
rect 317748 69136 317754 69148
rect 323578 69136 323584 69148
rect 317748 69108 323584 69136
rect 317748 69096 317754 69108
rect 323578 69096 323584 69108
rect 323636 69096 323642 69148
rect 345014 69096 345020 69148
rect 345072 69136 345078 69148
rect 349798 69136 349804 69148
rect 345072 69108 349804 69136
rect 345072 69096 345078 69108
rect 349798 69096 349804 69108
rect 349856 69096 349862 69148
rect 356606 69096 356612 69148
rect 356664 69136 356670 69148
rect 360838 69136 360844 69148
rect 356664 69108 360844 69136
rect 356664 69096 356670 69108
rect 360838 69096 360844 69108
rect 360896 69096 360902 69148
rect 104158 69028 104164 69080
rect 104216 69068 104222 69080
rect 104894 69068 104900 69080
rect 104216 69040 104900 69068
rect 104216 69028 104222 69040
rect 104894 69028 104900 69040
rect 104952 69028 104958 69080
rect 117958 69028 117964 69080
rect 118016 69068 118022 69080
rect 120534 69068 120540 69080
rect 118016 69040 120540 69068
rect 118016 69028 118022 69040
rect 120534 69028 120540 69040
rect 120592 69028 120598 69080
rect 162118 69028 162124 69080
rect 162176 69068 162182 69080
rect 165246 69068 165252 69080
rect 162176 69040 165252 69068
rect 162176 69028 162182 69040
rect 165246 69028 165252 69040
rect 165304 69028 165310 69080
rect 210418 69028 210424 69080
rect 210476 69068 210482 69080
rect 212534 69068 212540 69080
rect 210476 69040 212540 69068
rect 210476 69028 210482 69040
rect 212534 69028 212540 69040
rect 212592 69028 212598 69080
rect 224218 69028 224224 69080
rect 224276 69068 224282 69080
rect 224954 69068 224960 69080
rect 224276 69040 224960 69068
rect 224276 69028 224282 69040
rect 224954 69028 224960 69040
rect 225012 69028 225018 69080
rect 229738 69028 229744 69080
rect 229796 69068 229802 69080
rect 234798 69068 234804 69080
rect 229796 69040 234804 69068
rect 229796 69028 229802 69040
rect 234798 69028 234804 69040
rect 234856 69028 234862 69080
rect 242158 69028 242164 69080
rect 242216 69068 242222 69080
rect 243906 69068 243912 69080
rect 242216 69040 243912 69068
rect 242216 69028 242222 69040
rect 243906 69028 243912 69040
rect 243964 69028 243970 69080
rect 269758 69028 269764 69080
rect 269816 69068 269822 69080
rect 272058 69068 272064 69080
rect 269816 69040 272064 69068
rect 269816 69028 269822 69040
rect 272058 69028 272064 69040
rect 272116 69028 272122 69080
rect 279418 69028 279424 69080
rect 279476 69068 279482 69080
rect 281994 69068 282000 69080
rect 279476 69040 282000 69068
rect 279476 69028 279482 69040
rect 281994 69028 282000 69040
rect 282052 69028 282058 69080
rect 288434 69028 288440 69080
rect 288492 69068 288498 69080
rect 290274 69068 290280 69080
rect 288492 69040 290280 69068
rect 288492 69028 288498 69040
rect 290274 69028 290280 69040
rect 290332 69028 290338 69080
rect 298646 69028 298652 69080
rect 298704 69068 298710 69080
rect 299750 69068 299756 69080
rect 298704 69040 299756 69068
rect 298704 69028 298710 69040
rect 299750 69028 299756 69040
rect 299808 69028 299814 69080
rect 300302 69028 300308 69080
rect 300360 69068 300366 69080
rect 302234 69068 302240 69080
rect 300360 69040 302240 69068
rect 300360 69028 300366 69040
rect 302234 69028 302240 69040
rect 302292 69028 302298 69080
rect 304442 69028 304448 69080
rect 304500 69068 304506 69080
rect 305638 69068 305644 69080
rect 304500 69040 305644 69068
rect 304500 69028 304506 69040
rect 305638 69028 305644 69040
rect 305696 69028 305702 69080
rect 307754 69028 307760 69080
rect 307812 69068 307818 69080
rect 309778 69068 309784 69080
rect 307812 69040 309784 69068
rect 307812 69028 307818 69040
rect 309778 69028 309784 69040
rect 309836 69028 309842 69080
rect 312722 69028 312728 69080
rect 312780 69068 312786 69080
rect 313918 69068 313924 69080
rect 312780 69040 313924 69068
rect 312780 69028 312786 69040
rect 313918 69028 313924 69040
rect 313976 69028 313982 69080
rect 316034 69028 316040 69080
rect 316092 69068 316098 69080
rect 318058 69068 318064 69080
rect 316092 69040 318064 69068
rect 316092 69028 316098 69040
rect 318058 69028 318064 69040
rect 318116 69028 318122 69080
rect 330938 69028 330944 69080
rect 330996 69068 331002 69080
rect 331858 69068 331864 69080
rect 330996 69040 331864 69068
rect 330996 69028 331002 69040
rect 331858 69028 331864 69040
rect 331916 69028 331922 69080
rect 348326 69028 348332 69080
rect 348384 69068 348390 69080
rect 351178 69068 351184 69080
rect 348384 69040 351184 69068
rect 348384 69028 348390 69040
rect 351178 69028 351184 69040
rect 351236 69028 351242 69080
rect 355778 69028 355784 69080
rect 355836 69068 355842 69080
rect 356698 69068 356704 69080
rect 355836 69040 356704 69068
rect 355836 69028 355842 69040
rect 356698 69028 356704 69040
rect 356756 69028 356762 69080
rect 357434 69028 357440 69080
rect 357492 69068 357498 69080
rect 359458 69068 359464 69080
rect 357492 69040 359464 69068
rect 357492 69028 357498 69040
rect 359458 69028 359464 69040
rect 359516 69028 359522 69080
rect 362402 69028 362408 69080
rect 362460 69068 362466 69080
rect 363598 69068 363604 69080
rect 362460 69040 363604 69068
rect 362460 69028 362466 69040
rect 363598 69028 363604 69040
rect 363656 69028 363662 69080
rect 366542 69028 366548 69080
rect 366600 69068 366606 69080
rect 369118 69068 369124 69080
rect 366600 69040 369124 69068
rect 366600 69028 366606 69040
rect 369118 69028 369124 69040
rect 369176 69028 369182 69080
rect 398006 69028 398012 69080
rect 398064 69068 398070 69080
rect 399478 69068 399484 69080
rect 398064 69040 399484 69068
rect 398064 69028 398070 69040
rect 399478 69028 399484 69040
rect 399536 69028 399542 69080
rect 438578 69028 438584 69080
rect 438636 69068 438642 69080
rect 439498 69068 439504 69080
rect 438636 69040 439504 69068
rect 438636 69028 438642 69040
rect 439498 69028 439504 69040
rect 439556 69028 439562 69080
rect 443546 69028 443552 69080
rect 443604 69068 443610 69080
rect 445018 69068 445024 69080
rect 443604 69040 445024 69068
rect 443604 69028 443610 69040
rect 445018 69028 445024 69040
rect 445076 69028 445082 69080
rect 455966 69028 455972 69080
rect 456024 69068 456030 69080
rect 458818 69068 458824 69080
rect 456024 69040 458824 69068
rect 456024 69028 456030 69040
rect 458818 69028 458824 69040
rect 458876 69028 458882 69080
rect 460934 69028 460940 69080
rect 460992 69068 460998 69080
rect 468478 69068 468484 69080
rect 460992 69040 468484 69068
rect 460992 69028 460998 69040
rect 468478 69028 468484 69040
rect 468536 69028 468542 69080
rect 470870 69028 470876 69080
rect 470928 69068 470934 69080
rect 472618 69068 472624 69080
rect 470928 69040 472624 69068
rect 470928 69028 470934 69040
rect 472618 69028 472624 69040
rect 472676 69028 472682 69080
rect 475838 69028 475844 69080
rect 475896 69068 475902 69080
rect 476758 69068 476764 69080
rect 475896 69040 476764 69068
rect 475896 69028 475902 69040
rect 476758 69028 476764 69040
rect 476816 69028 476822 69080
rect 480806 69028 480812 69080
rect 480864 69068 480870 69080
rect 482278 69068 482284 69080
rect 480864 69040 482284 69068
rect 480864 69028 480870 69040
rect 482278 69028 482284 69040
rect 482336 69028 482342 69080
rect 207014 68416 207020 68468
rect 207072 68456 207078 68468
rect 233234 68456 233240 68468
rect 207072 68428 233240 68456
rect 207072 68416 207078 68428
rect 233234 68416 233240 68428
rect 233292 68416 233298 68468
rect 253198 68416 253204 68468
rect 253256 68456 253262 68468
rect 256326 68456 256332 68468
rect 253256 68428 256332 68456
rect 253256 68416 253262 68428
rect 256326 68416 256332 68428
rect 256384 68416 256390 68468
rect 149054 68348 149060 68400
rect 149112 68388 149118 68400
rect 192570 68388 192576 68400
rect 149112 68360 192576 68388
rect 149112 68348 149118 68360
rect 192570 68348 192576 68360
rect 192628 68348 192634 68400
rect 193214 68348 193220 68400
rect 193272 68388 193278 68400
rect 223206 68388 223212 68400
rect 193272 68360 223212 68388
rect 193272 68348 193278 68360
rect 223206 68348 223212 68360
rect 223264 68348 223270 68400
rect 370682 68348 370688 68400
rect 370740 68388 370746 68400
rect 402974 68388 402980 68400
rect 370740 68360 402980 68388
rect 370740 68348 370746 68360
rect 402974 68348 402980 68360
rect 403032 68348 403038 68400
rect 434438 68348 434444 68400
rect 434496 68388 434502 68400
rect 494146 68388 494152 68400
rect 434496 68360 494152 68388
rect 434496 68348 434502 68360
rect 494146 68348 494152 68360
rect 494204 68348 494210 68400
rect 7558 68280 7564 68332
rect 7616 68320 7622 68332
rect 89070 68320 89076 68332
rect 7616 68292 89076 68320
rect 7616 68280 7622 68292
rect 89070 68280 89076 68292
rect 89128 68280 89134 68332
rect 93854 68280 93860 68332
rect 93912 68320 93918 68332
rect 154574 68320 154580 68332
rect 93912 68292 154580 68320
rect 93912 68280 93918 68292
rect 154574 68280 154580 68292
rect 154632 68280 154638 68332
rect 171134 68280 171140 68332
rect 171192 68320 171198 68332
rect 208394 68320 208400 68332
rect 171192 68292 208400 68320
rect 171192 68280 171198 68292
rect 208394 68280 208400 68292
rect 208452 68280 208458 68332
rect 227714 68280 227720 68332
rect 227772 68320 227778 68332
rect 248046 68320 248052 68332
rect 227772 68292 248052 68320
rect 227772 68280 227778 68292
rect 248046 68280 248052 68292
rect 248104 68280 248110 68332
rect 249794 68280 249800 68332
rect 249852 68320 249858 68332
rect 262950 68320 262956 68332
rect 249852 68292 262956 68320
rect 249852 68280 249858 68292
rect 262950 68280 262956 68292
rect 263008 68280 263014 68332
rect 383930 68280 383936 68332
rect 383988 68320 383994 68332
rect 422294 68320 422300 68332
rect 383988 68292 422300 68320
rect 383988 68280 383994 68292
rect 422294 68280 422300 68292
rect 422352 68280 422358 68332
rect 465074 68280 465080 68332
rect 465132 68320 465138 68332
rect 538214 68320 538220 68332
rect 465132 68292 538220 68320
rect 465132 68280 465138 68292
rect 538214 68280 538220 68292
rect 538272 68280 538278 68332
rect 489914 67600 489920 67652
rect 489972 67640 489978 67652
rect 490190 67640 490196 67652
rect 489972 67612 490196 67640
rect 489972 67600 489978 67612
rect 490190 67600 490196 67612
rect 490248 67600 490254 67652
rect 209774 67056 209780 67108
rect 209832 67096 209838 67108
rect 235626 67096 235632 67108
rect 209832 67068 235632 67096
rect 209832 67056 209838 67068
rect 235626 67056 235632 67068
rect 235684 67056 235690 67108
rect 200114 66988 200120 67040
rect 200172 67028 200178 67040
rect 228174 67028 228180 67040
rect 200172 67000 228180 67028
rect 200172 66988 200178 67000
rect 228174 66988 228180 67000
rect 228232 66988 228238 67040
rect 80054 66920 80060 66972
rect 80112 66960 80118 66972
rect 144546 66960 144552 66972
rect 80112 66932 144552 66960
rect 80112 66920 80118 66932
rect 144546 66920 144552 66932
rect 144604 66920 144610 66972
rect 165614 66920 165620 66972
rect 165672 66960 165678 66972
rect 204254 66960 204260 66972
rect 165672 66932 204260 66960
rect 165672 66920 165678 66932
rect 204254 66920 204260 66932
rect 204312 66920 204318 66972
rect 4798 66852 4804 66904
rect 4856 66892 4862 66904
rect 88334 66892 88340 66904
rect 4856 66864 88340 66892
rect 4856 66852 4862 66864
rect 88334 66852 88340 66864
rect 88392 66852 88398 66904
rect 115934 66852 115940 66904
rect 115992 66892 115998 66904
rect 169386 66892 169392 66904
rect 115992 66864 169392 66892
rect 115992 66852 115998 66864
rect 169386 66852 169392 66864
rect 169444 66852 169450 66904
rect 175274 66852 175280 66904
rect 175332 66892 175338 66904
rect 210786 66892 210792 66904
rect 175332 66864 210792 66892
rect 175332 66852 175338 66864
rect 210786 66852 210792 66864
rect 210844 66852 210850 66904
rect 238754 66852 238760 66904
rect 238812 66892 238818 66904
rect 255498 66892 255504 66904
rect 238812 66864 255504 66892
rect 238812 66852 238818 66864
rect 255498 66852 255504 66864
rect 255556 66852 255562 66904
rect 375650 66852 375656 66904
rect 375708 66892 375714 66904
rect 409874 66892 409880 66904
rect 375708 66864 409880 66892
rect 375708 66852 375714 66864
rect 409874 66852 409880 66864
rect 409932 66852 409938 66904
rect 479150 66852 479156 66904
rect 479208 66892 479214 66904
rect 557534 66892 557540 66904
rect 479208 66864 557540 66892
rect 479208 66852 479214 66864
rect 557534 66852 557540 66864
rect 557592 66852 557598 66904
rect 255958 66240 255964 66292
rect 256016 66280 256022 66292
rect 259638 66280 259644 66292
rect 256016 66252 259644 66280
rect 256016 66240 256022 66252
rect 259638 66240 259644 66252
rect 259696 66240 259702 66292
rect 324406 66172 324412 66224
rect 324464 66212 324470 66224
rect 325050 66212 325056 66224
rect 324464 66184 325056 66212
rect 324464 66172 324470 66184
rect 325050 66172 325056 66184
rect 325108 66172 325114 66224
rect 224954 65764 224960 65816
rect 225012 65804 225018 65816
rect 245654 65804 245660 65816
rect 225012 65776 245660 65804
rect 225012 65764 225018 65776
rect 245654 65764 245660 65776
rect 245712 65764 245718 65816
rect 196066 65628 196072 65680
rect 196124 65668 196130 65680
rect 225690 65668 225696 65680
rect 196124 65640 225696 65668
rect 196124 65628 196130 65640
rect 225690 65628 225696 65640
rect 225748 65628 225754 65680
rect 259546 65628 259552 65680
rect 259604 65668 259610 65680
rect 269574 65668 269580 65680
rect 259604 65640 269580 65668
rect 259604 65628 259610 65640
rect 269574 65628 269580 65640
rect 269632 65628 269638 65680
rect 44174 65492 44180 65544
rect 44232 65532 44238 65544
rect 118878 65532 118884 65544
rect 44232 65504 118884 65532
rect 44232 65492 44238 65504
rect 118878 65492 118884 65504
rect 118936 65492 118942 65544
rect 157978 65492 157984 65544
rect 158036 65532 158042 65544
rect 196710 65532 196716 65544
rect 158036 65504 196716 65532
rect 158036 65492 158042 65504
rect 196710 65492 196716 65504
rect 196768 65492 196774 65544
rect 211154 65492 211160 65544
rect 211212 65532 211218 65544
rect 236454 65532 236460 65544
rect 211212 65504 236460 65532
rect 211212 65492 211218 65504
rect 236454 65492 236460 65504
rect 236512 65492 236518 65544
rect 245654 65492 245660 65544
rect 245712 65532 245718 65544
rect 260466 65532 260472 65544
rect 245712 65504 260472 65532
rect 245712 65492 245718 65504
rect 260466 65492 260472 65504
rect 260524 65492 260530 65544
rect 402146 65492 402152 65544
rect 402204 65532 402210 65544
rect 448514 65532 448520 65544
rect 402204 65504 448520 65532
rect 402204 65492 402210 65504
rect 448514 65492 448520 65504
rect 448572 65492 448578 65544
rect 484118 65492 484124 65544
rect 484176 65532 484182 65544
rect 564526 65532 564532 65544
rect 484176 65504 564532 65532
rect 484176 65492 484182 65504
rect 564526 65492 564532 65504
rect 564584 65492 564590 65544
rect 146386 64336 146392 64388
rect 146444 64376 146450 64388
rect 190454 64376 190460 64388
rect 146444 64348 190460 64376
rect 146444 64336 146450 64348
rect 190454 64336 190460 64348
rect 190512 64336 190518 64388
rect 220814 64336 220820 64388
rect 220872 64376 220878 64388
rect 242986 64376 242992 64388
rect 220872 64348 242992 64376
rect 220872 64336 220878 64348
rect 242986 64336 242992 64348
rect 243044 64336 243050 64388
rect 84194 64200 84200 64252
rect 84252 64240 84258 64252
rect 146478 64240 146484 64252
rect 84252 64212 146484 64240
rect 84252 64200 84258 64212
rect 146478 64200 146484 64212
rect 146536 64200 146542 64252
rect 192478 64200 192484 64252
rect 192536 64240 192542 64252
rect 220998 64240 221004 64252
rect 192536 64212 221004 64240
rect 192536 64200 192542 64212
rect 220998 64200 221004 64212
rect 221056 64200 221062 64252
rect 28994 64132 29000 64184
rect 29052 64172 29058 64184
rect 109034 64172 109040 64184
rect 29052 64144 109040 64172
rect 29052 64132 29058 64144
rect 109034 64132 109040 64144
rect 109092 64132 109098 64184
rect 189166 64132 189172 64184
rect 189224 64172 189230 64184
rect 220906 64172 220912 64184
rect 189224 64144 220912 64172
rect 189224 64132 189230 64144
rect 220906 64132 220912 64144
rect 220964 64132 220970 64184
rect 242986 64132 242992 64184
rect 243044 64172 243050 64184
rect 258074 64172 258080 64184
rect 243044 64144 258080 64172
rect 243044 64132 243050 64144
rect 258074 64132 258080 64144
rect 258132 64132 258138 64184
rect 481634 64132 481640 64184
rect 481692 64172 481698 64184
rect 561674 64172 561680 64184
rect 481692 64144 561680 64172
rect 481692 64132 481698 64144
rect 561674 64132 561680 64144
rect 561732 64132 561738 64184
rect 121546 62908 121552 62960
rect 121604 62948 121610 62960
rect 172606 62948 172612 62960
rect 121604 62920 172612 62948
rect 121604 62908 121610 62920
rect 172606 62908 172612 62920
rect 172664 62908 172670 62960
rect 444374 62840 444380 62892
rect 444432 62880 444438 62892
rect 507854 62880 507860 62892
rect 444432 62852 507860 62880
rect 444432 62840 444438 62852
rect 507854 62840 507860 62852
rect 507912 62840 507918 62892
rect 46934 62772 46940 62824
rect 46992 62812 46998 62824
rect 121638 62812 121644 62824
rect 46992 62784 121644 62812
rect 46992 62772 46998 62784
rect 121638 62772 121644 62784
rect 121696 62772 121702 62824
rect 178034 62772 178040 62824
rect 178092 62812 178098 62824
rect 212626 62812 212632 62824
rect 178092 62784 212632 62812
rect 178092 62772 178098 62784
rect 212626 62772 212632 62784
rect 212684 62772 212690 62824
rect 214006 62772 214012 62824
rect 214064 62812 214070 62824
rect 237466 62812 237472 62824
rect 214064 62784 237472 62812
rect 214064 62772 214070 62784
rect 237466 62772 237472 62784
rect 237524 62772 237530 62824
rect 478874 62772 478880 62824
rect 478932 62812 478938 62824
rect 558914 62812 558920 62824
rect 478932 62784 558920 62812
rect 478932 62772 478938 62784
rect 558914 62772 558920 62784
rect 558972 62772 558978 62824
rect 484394 61344 484400 61396
rect 484452 61384 484458 61396
rect 565814 61384 565820 61396
rect 484452 61356 565820 61384
rect 484452 61344 484458 61356
rect 565814 61344 565820 61356
rect 565872 61344 565878 61396
rect 577866 60664 577872 60716
rect 577924 60704 577930 60716
rect 579982 60704 579988 60716
rect 577924 60676 579988 60704
rect 577924 60664 577930 60676
rect 579982 60664 579988 60676
rect 580040 60664 580046 60716
rect 13078 59984 13084 60036
rect 13136 60024 13142 60036
rect 94222 60024 94228 60036
rect 13136 59996 94228 60024
rect 13136 59984 13142 59996
rect 94222 59984 94228 59996
rect 94280 59984 94286 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 512086 59344 512092 59356
rect 3108 59316 512092 59344
rect 3108 59304 3114 59316
rect 512086 59304 512092 59316
rect 512144 59304 512150 59356
rect 74534 58692 74540 58744
rect 74592 58732 74598 58744
rect 139486 58732 139492 58744
rect 74592 58704 139492 58732
rect 74592 58692 74598 58704
rect 139486 58692 139492 58704
rect 139544 58692 139550 58744
rect 27614 58624 27620 58676
rect 27672 58664 27678 58676
rect 106642 58664 106648 58676
rect 27672 58636 106648 58664
rect 27672 58624 27678 58636
rect 106642 58624 106648 58636
rect 106700 58624 106706 58676
rect 174630 58624 174636 58676
rect 174688 58664 174694 58676
rect 208578 58664 208584 58676
rect 174688 58636 208584 58664
rect 174688 58624 174694 58636
rect 208578 58624 208584 58636
rect 208636 58624 208642 58676
rect 469306 58624 469312 58676
rect 469364 58664 469370 58676
rect 545114 58664 545120 58676
rect 469364 58636 545120 58664
rect 469364 58624 469370 58636
rect 545114 58624 545120 58636
rect 545172 58624 545178 58676
rect 67634 57264 67640 57316
rect 67692 57304 67698 57316
rect 135346 57304 135352 57316
rect 67692 57276 135352 57304
rect 67692 57264 67698 57276
rect 135346 57264 135352 57276
rect 135404 57264 135410 57316
rect 429286 57264 429292 57316
rect 429344 57304 429350 57316
rect 488626 57304 488632 57316
rect 429344 57276 488632 57304
rect 429344 57264 429350 57276
rect 488626 57264 488632 57276
rect 488684 57264 488690 57316
rect 17954 57196 17960 57248
rect 18012 57236 18018 57248
rect 100754 57236 100760 57248
rect 18012 57208 100760 57236
rect 18012 57196 18018 57208
rect 100754 57196 100760 57208
rect 100812 57196 100818 57248
rect 182818 57196 182824 57248
rect 182876 57236 182882 57248
rect 214098 57236 214104 57248
rect 182876 57208 214104 57236
rect 182876 57196 182882 57208
rect 214098 57196 214104 57208
rect 214156 57196 214162 57248
rect 473354 57196 473360 57248
rect 473412 57236 473418 57248
rect 549254 57236 549260 57248
rect 473412 57208 549260 57236
rect 473412 57196 473418 57208
rect 549254 57196 549260 57208
rect 549312 57196 549318 57248
rect 30374 55836 30380 55888
rect 30432 55876 30438 55888
rect 109218 55876 109224 55888
rect 30432 55848 109224 55876
rect 30432 55836 30438 55848
rect 109218 55836 109224 55848
rect 109276 55836 109282 55888
rect 144914 55836 144920 55888
rect 144972 55876 144978 55888
rect 189442 55876 189448 55888
rect 144972 55848 189448 55876
rect 144972 55836 144978 55848
rect 189442 55836 189448 55848
rect 189500 55836 189506 55888
rect 415394 55836 415400 55888
rect 415452 55876 415458 55888
rect 466546 55876 466552 55888
rect 415452 55848 466552 55876
rect 415452 55836 415458 55848
rect 466546 55836 466552 55848
rect 466604 55836 466610 55888
rect 487154 55836 487160 55888
rect 487212 55876 487218 55888
rect 569954 55876 569960 55888
rect 487212 55848 569960 55876
rect 487212 55836 487218 55848
rect 569954 55836 569960 55848
rect 570012 55836 570018 55888
rect 433334 54544 433340 54596
rect 433392 54584 433398 54596
rect 492674 54584 492680 54596
rect 433392 54556 492680 54584
rect 433392 54544 433398 54556
rect 492674 54544 492680 54556
rect 492732 54544 492738 54596
rect 44266 54476 44272 54528
rect 44324 54516 44330 54528
rect 118694 54516 118700 54528
rect 44324 54488 118700 54516
rect 44324 54476 44330 54488
rect 118694 54476 118700 54488
rect 118752 54476 118758 54528
rect 490006 54476 490012 54528
rect 490064 54516 490070 54528
rect 574094 54516 574100 54528
rect 490064 54488 574100 54516
rect 490064 54476 490070 54488
rect 574094 54476 574100 54488
rect 574152 54476 574158 54528
rect 41414 53048 41420 53100
rect 41472 53088 41478 53100
rect 117314 53088 117320 53100
rect 41472 53060 117320 53088
rect 41472 53048 41478 53060
rect 117314 53048 117320 53060
rect 117372 53048 117378 53100
rect 491386 53048 491392 53100
rect 491444 53088 491450 53100
rect 576118 53088 576124 53100
rect 491444 53060 576124 53088
rect 491444 53048 491450 53060
rect 576118 53048 576124 53060
rect 576176 53048 576182 53100
rect 37274 51688 37280 51740
rect 37332 51728 37338 51740
rect 114646 51728 114652 51740
rect 37332 51700 114652 51728
rect 37332 51688 37338 51700
rect 114646 51688 114652 51700
rect 114704 51688 114710 51740
rect 151814 51688 151820 51740
rect 151872 51728 151878 51740
rect 194594 51728 194600 51740
rect 151872 51700 194600 51728
rect 151872 51688 151878 51700
rect 194594 51688 194600 51700
rect 194652 51688 194658 51740
rect 440326 51688 440332 51740
rect 440384 51728 440390 51740
rect 503714 51728 503720 51740
rect 440384 51700 503720 51728
rect 440384 51688 440390 51700
rect 503714 51688 503720 51700
rect 503772 51688 503778 51740
rect 102226 50396 102232 50448
rect 102284 50436 102290 50448
rect 158806 50436 158812 50448
rect 102284 50408 158812 50436
rect 102284 50396 102290 50408
rect 158806 50396 158812 50408
rect 158864 50396 158870 50448
rect 24854 50328 24860 50380
rect 24912 50368 24918 50380
rect 104986 50368 104992 50380
rect 24912 50340 104992 50368
rect 24912 50328 24918 50340
rect 104986 50328 104992 50340
rect 105044 50328 105050 50380
rect 188338 50328 188344 50380
rect 188396 50368 188402 50380
rect 218146 50368 218152 50380
rect 188396 50340 218152 50368
rect 188396 50328 188402 50340
rect 218146 50328 218152 50340
rect 218204 50328 218210 50380
rect 439498 50328 439504 50380
rect 439556 50368 439562 50380
rect 499574 50368 499580 50380
rect 439556 50340 499580 50368
rect 439556 50328 439562 50340
rect 499574 50328 499580 50340
rect 499632 50328 499638 50380
rect 92658 49036 92664 49088
rect 92716 49076 92722 49088
rect 152182 49076 152188 49088
rect 92716 49048 152188 49076
rect 92716 49036 92722 49048
rect 152182 49036 152188 49048
rect 152240 49036 152246 49088
rect 425146 49036 425152 49088
rect 425204 49076 425210 49088
rect 481634 49076 481640 49088
rect 425204 49048 481640 49076
rect 425204 49036 425210 49048
rect 481634 49036 481640 49048
rect 481692 49036 481698 49088
rect 49694 48968 49700 49020
rect 49752 49008 49758 49020
rect 122926 49008 122932 49020
rect 49752 48980 122932 49008
rect 49752 48968 49758 48980
rect 122926 48968 122932 48980
rect 122984 48968 122990 49020
rect 218146 48968 218152 49020
rect 218204 49008 218210 49020
rect 240134 49008 240140 49020
rect 218204 48980 240140 49008
rect 218204 48968 218210 48980
rect 240134 48968 240140 48980
rect 240192 48968 240198 49020
rect 449986 48968 449992 49020
rect 450044 49008 450050 49020
rect 517514 49008 517520 49020
rect 450044 48980 517520 49008
rect 450044 48968 450050 48980
rect 517514 48968 517520 48980
rect 517572 48968 517578 49020
rect 512638 46860 512644 46912
rect 512696 46900 512702 46912
rect 580166 46900 580172 46912
rect 512696 46872 580172 46900
rect 512696 46860 512702 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 60734 46180 60740 46232
rect 60792 46220 60798 46232
rect 131206 46220 131212 46232
rect 60792 46192 131212 46220
rect 60792 46180 60798 46192
rect 131206 46180 131212 46192
rect 131264 46180 131270 46232
rect 400214 46180 400220 46232
rect 400272 46220 400278 46232
rect 445754 46220 445760 46232
rect 400272 46192 445760 46220
rect 400272 46180 400278 46192
rect 445754 46180 445760 46192
rect 445812 46180 445818 46232
rect 445846 46180 445852 46232
rect 445904 46220 445910 46232
rect 512086 46220 512092 46232
rect 445904 46192 512092 46220
rect 445904 46180 445910 46192
rect 512086 46180 512092 46192
rect 512144 46180 512150 46232
rect 110506 44888 110512 44940
rect 110564 44928 110570 44940
rect 162118 44928 162124 44940
rect 110564 44900 162124 44928
rect 110564 44888 110570 44900
rect 162118 44888 162124 44900
rect 162176 44888 162182 44940
rect 431954 44888 431960 44940
rect 432012 44928 432018 44940
rect 489914 44928 489920 44940
rect 432012 44900 489920 44928
rect 432012 44888 432018 44900
rect 489914 44888 489920 44900
rect 489972 44888 489978 44940
rect 53834 44820 53840 44872
rect 53892 44860 53898 44872
rect 125686 44860 125692 44872
rect 53892 44832 125692 44860
rect 53892 44820 53898 44832
rect 125686 44820 125692 44832
rect 125744 44820 125750 44872
rect 223666 44820 223672 44872
rect 223724 44860 223730 44872
rect 244274 44860 244280 44872
rect 223724 44832 244280 44860
rect 223724 44820 223730 44832
rect 244274 44820 244280 44832
rect 244332 44820 244338 44872
rect 379606 44820 379612 44872
rect 379664 44860 379670 44872
rect 416866 44860 416872 44872
rect 379664 44832 416872 44860
rect 379664 44820 379670 44832
rect 416866 44820 416872 44832
rect 416924 44820 416930 44872
rect 458818 44820 458824 44872
rect 458876 44860 458882 44872
rect 524414 44860 524420 44872
rect 458876 44832 524420 44860
rect 458876 44820 458882 44832
rect 524414 44820 524420 44832
rect 524472 44820 524478 44872
rect 63494 43460 63500 43512
rect 63552 43500 63558 43512
rect 132494 43500 132500 43512
rect 63552 43472 132500 43500
rect 63552 43460 63558 43472
rect 132494 43460 132500 43472
rect 132552 43460 132558 43512
rect 436094 43460 436100 43512
rect 436152 43500 436158 43512
rect 496814 43500 496820 43512
rect 436152 43472 496820 43500
rect 436152 43460 436158 43472
rect 496814 43460 496820 43472
rect 496872 43460 496878 43512
rect 17218 43392 17224 43444
rect 17276 43432 17282 43444
rect 96706 43432 96712 43444
rect 17276 43404 96712 43432
rect 17276 43392 17282 43404
rect 96706 43392 96712 43404
rect 96764 43392 96770 43444
rect 142246 43392 142252 43444
rect 142304 43432 142310 43444
rect 187694 43432 187700 43444
rect 142304 43404 187700 43432
rect 142304 43392 142310 43404
rect 187694 43392 187700 43404
rect 187752 43392 187758 43444
rect 476758 43392 476764 43444
rect 476816 43432 476822 43444
rect 553394 43432 553400 43444
rect 476816 43404 553400 43432
rect 476816 43392 476822 43404
rect 553394 43392 553400 43404
rect 553452 43392 553458 43444
rect 56594 42100 56600 42152
rect 56652 42140 56658 42152
rect 127066 42140 127072 42152
rect 56652 42112 127072 42140
rect 56652 42100 56658 42112
rect 127066 42100 127072 42112
rect 127124 42100 127130 42152
rect 8938 42032 8944 42084
rect 8996 42072 9002 42084
rect 89806 42072 89812 42084
rect 8996 42044 89812 42072
rect 8996 42032 9002 42044
rect 89806 42032 89812 42044
rect 89864 42032 89870 42084
rect 102318 42032 102324 42084
rect 102376 42072 102382 42084
rect 160186 42072 160192 42084
rect 102376 42044 160192 42072
rect 102376 42032 102382 42044
rect 160186 42032 160192 42044
rect 160244 42032 160250 42084
rect 231854 42032 231860 42084
rect 231912 42072 231918 42084
rect 249886 42072 249892 42084
rect 231912 42044 249892 42072
rect 231912 42032 231918 42044
rect 249886 42032 249892 42044
rect 249944 42032 249950 42084
rect 419626 42032 419632 42084
rect 419684 42072 419690 42084
rect 473354 42072 473360 42084
rect 419684 42044 473360 42072
rect 419684 42032 419690 42044
rect 473354 42032 473360 42044
rect 473412 42032 473418 42084
rect 481726 42032 481732 42084
rect 481784 42072 481790 42084
rect 563054 42072 563060 42084
rect 481784 42044 563060 42072
rect 481784 42032 481790 42044
rect 563054 42032 563060 42044
rect 563112 42032 563118 42084
rect 99466 40740 99472 40792
rect 99524 40780 99530 40792
rect 157334 40780 157340 40792
rect 99524 40752 157340 40780
rect 99524 40740 99530 40752
rect 157334 40740 157340 40752
rect 157392 40740 157398 40792
rect 52454 40672 52460 40724
rect 52512 40712 52518 40724
rect 125594 40712 125600 40724
rect 52512 40684 125600 40712
rect 52512 40672 52518 40684
rect 125594 40672 125600 40684
rect 125652 40672 125658 40724
rect 436186 40672 436192 40724
rect 436244 40712 436250 40724
rect 498194 40712 498200 40724
rect 436244 40684 498200 40712
rect 436244 40672 436250 40684
rect 498194 40672 498200 40684
rect 498252 40672 498258 40724
rect 111794 39448 111800 39500
rect 111852 39488 111858 39500
rect 166994 39488 167000 39500
rect 111852 39460 167000 39488
rect 111852 39448 111858 39460
rect 166994 39448 167000 39460
rect 167052 39448 167058 39500
rect 423674 39380 423680 39432
rect 423732 39420 423738 39432
rect 478874 39420 478880 39432
rect 423732 39392 478880 39420
rect 423732 39380 423738 39392
rect 478874 39380 478880 39392
rect 478932 39380 478938 39432
rect 34514 39312 34520 39364
rect 34572 39352 34578 39364
rect 111886 39352 111892 39364
rect 34572 39324 111892 39352
rect 34572 39312 34578 39324
rect 111886 39312 111892 39324
rect 111944 39312 111950 39364
rect 477494 39312 477500 39364
rect 477552 39352 477558 39364
rect 556246 39352 556252 39364
rect 477552 39324 556252 39352
rect 477552 39312 477558 39324
rect 556246 39312 556252 39324
rect 556304 39312 556310 39364
rect 85574 37952 85580 38004
rect 85632 37992 85638 38004
rect 147766 37992 147772 38004
rect 85632 37964 147772 37992
rect 85632 37952 85638 37964
rect 147766 37952 147772 37964
rect 147824 37952 147830 38004
rect 432046 37952 432052 38004
rect 432104 37992 432110 38004
rect 491386 37992 491392 38004
rect 432104 37964 491392 37992
rect 432104 37952 432110 37964
rect 491386 37952 491392 37964
rect 491444 37952 491450 38004
rect 35894 37884 35900 37936
rect 35952 37924 35958 37936
rect 113266 37924 113272 37936
rect 35952 37896 113272 37924
rect 35952 37884 35958 37896
rect 113266 37884 113272 37896
rect 113324 37884 113330 37936
rect 485774 37884 485780 37936
rect 485832 37924 485838 37936
rect 567194 37924 567200 37936
rect 485832 37896 567200 37924
rect 485832 37884 485838 37896
rect 567194 37884 567200 37896
rect 567252 37884 567258 37936
rect 26234 36524 26240 36576
rect 26292 36564 26298 36576
rect 106366 36564 106372 36576
rect 26292 36536 106372 36564
rect 26292 36524 26298 36536
rect 106366 36524 106372 36536
rect 106424 36524 106430 36576
rect 118694 36524 118700 36576
rect 118752 36564 118758 36576
rect 171318 36564 171324 36576
rect 118752 36536 171324 36564
rect 118752 36524 118758 36536
rect 171318 36524 171324 36536
rect 171376 36524 171382 36576
rect 445018 36524 445024 36576
rect 445076 36564 445082 36576
rect 506474 36564 506480 36576
rect 445076 36536 506480 36564
rect 445076 36524 445082 36536
rect 506474 36524 506480 36536
rect 506532 36524 506538 36576
rect 98178 35164 98184 35216
rect 98236 35204 98242 35216
rect 156046 35204 156052 35216
rect 98236 35176 156052 35204
rect 98236 35164 98242 35176
rect 156046 35164 156052 35176
rect 156104 35164 156110 35216
rect 430574 35164 430580 35216
rect 430632 35204 430638 35216
rect 490006 35204 490012 35216
rect 430632 35176 490012 35204
rect 430632 35164 430638 35176
rect 490006 35164 490012 35176
rect 490064 35164 490070 35216
rect 31754 33736 31760 33788
rect 31812 33776 31818 33788
rect 110598 33776 110604 33788
rect 31812 33748 110604 33776
rect 31812 33736 31818 33748
rect 110598 33736 110604 33748
rect 110656 33736 110662 33788
rect 114646 33736 114652 33788
rect 114704 33776 114710 33788
rect 168374 33776 168380 33788
rect 114704 33748 168380 33776
rect 114704 33736 114710 33748
rect 168374 33736 168380 33748
rect 168432 33736 168438 33788
rect 427906 33736 427912 33788
rect 427964 33776 427970 33788
rect 485774 33776 485780 33788
rect 427964 33748 485780 33776
rect 427964 33736 427970 33748
rect 485774 33736 485780 33748
rect 485832 33736 485838 33788
rect 490190 33736 490196 33788
rect 490248 33776 490254 33788
rect 572714 33776 572720 33788
rect 490248 33748 572720 33776
rect 490248 33736 490254 33748
rect 572714 33736 572720 33748
rect 572772 33736 572778 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 72418 33096 72424 33108
rect 3200 33068 72424 33096
rect 3200 33056 3206 33068
rect 72418 33056 72424 33068
rect 72476 33056 72482 33108
rect 514018 33056 514024 33108
rect 514076 33096 514082 33108
rect 580166 33096 580172 33108
rect 514076 33068 580172 33096
rect 514076 33056 514082 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 417142 32444 417148 32496
rect 417200 32484 417206 32496
rect 470686 32484 470692 32496
rect 417200 32456 470692 32484
rect 417200 32444 417206 32456
rect 470686 32444 470692 32456
rect 470744 32444 470750 32496
rect 107654 32376 107660 32428
rect 107712 32416 107718 32428
rect 162946 32416 162952 32428
rect 107712 32388 162952 32416
rect 107712 32376 107718 32388
rect 162946 32376 162952 32388
rect 163004 32376 163010 32428
rect 453298 32376 453304 32428
rect 453356 32416 453362 32428
rect 510614 32416 510620 32428
rect 453356 32388 510620 32416
rect 453356 32376 453362 32388
rect 510614 32376 510620 32388
rect 510672 32376 510678 32428
rect 91094 31016 91100 31068
rect 91152 31056 91158 31068
rect 151906 31056 151912 31068
rect 91152 31028 151912 31056
rect 91152 31016 91158 31028
rect 151906 31016 151912 31028
rect 151964 31016 151970 31068
rect 156046 31016 156052 31068
rect 156104 31056 156110 31068
rect 197538 31056 197544 31068
rect 156104 31028 197544 31056
rect 156104 31016 156110 31028
rect 197538 31016 197544 31028
rect 197596 31016 197602 31068
rect 390554 31016 390560 31068
rect 390612 31056 390618 31068
rect 432046 31056 432052 31068
rect 390612 31028 432052 31056
rect 390612 31016 390618 31028
rect 432046 31016 432052 31028
rect 432104 31016 432110 31068
rect 454126 31016 454132 31068
rect 454184 31056 454190 31068
rect 523034 31056 523040 31068
rect 454184 31028 523040 31056
rect 454184 31016 454190 31028
rect 523034 31016 523040 31028
rect 523092 31016 523098 31068
rect 60826 29588 60832 29640
rect 60884 29628 60890 29640
rect 129826 29628 129832 29640
rect 60884 29600 129832 29628
rect 60884 29588 60890 29600
rect 129826 29588 129832 29600
rect 129884 29588 129890 29640
rect 135346 29588 135352 29640
rect 135404 29628 135410 29640
rect 182174 29628 182180 29640
rect 135404 29600 182180 29628
rect 135404 29588 135410 29600
rect 182174 29588 182180 29600
rect 182232 29588 182238 29640
rect 412726 29588 412732 29640
rect 412784 29628 412790 29640
rect 463786 29628 463792 29640
rect 412784 29600 463792 29628
rect 412784 29588 412790 29600
rect 463786 29588 463792 29600
rect 463844 29588 463850 29640
rect 471974 29588 471980 29640
rect 472032 29628 472038 29640
rect 547874 29628 547880 29640
rect 472032 29600 547880 29628
rect 472032 29588 472038 29600
rect 547874 29588 547880 29600
rect 547932 29588 547938 29640
rect 86954 28228 86960 28280
rect 87012 28268 87018 28280
rect 149146 28268 149152 28280
rect 87012 28240 149152 28268
rect 87012 28228 87018 28240
rect 149146 28228 149152 28240
rect 149204 28228 149210 28280
rect 151906 28228 151912 28280
rect 151964 28268 151970 28280
rect 193582 28268 193588 28280
rect 151964 28240 193588 28268
rect 151964 28228 151970 28240
rect 193582 28228 193588 28240
rect 193640 28228 193646 28280
rect 382366 28228 382372 28280
rect 382424 28268 382430 28280
rect 421006 28268 421012 28280
rect 382424 28240 421012 28268
rect 382424 28228 382430 28240
rect 421006 28228 421012 28240
rect 421064 28228 421070 28280
rect 425054 28228 425060 28280
rect 425112 28268 425118 28280
rect 481726 28268 481732 28280
rect 425112 28240 481732 28268
rect 425112 28228 425118 28240
rect 481726 28228 481732 28240
rect 481784 28228 481790 28280
rect 73154 26868 73160 26920
rect 73212 26908 73218 26920
rect 139394 26908 139400 26920
rect 73212 26880 139400 26908
rect 73212 26868 73218 26880
rect 139394 26868 139400 26880
rect 139452 26868 139458 26920
rect 147766 26868 147772 26920
rect 147824 26908 147830 26920
rect 191926 26908 191932 26920
rect 147824 26880 191932 26908
rect 147824 26868 147830 26880
rect 191926 26868 191932 26880
rect 191984 26868 191990 26920
rect 409966 26868 409972 26920
rect 410024 26908 410030 26920
rect 459646 26908 459652 26920
rect 410024 26880 459652 26908
rect 410024 26868 410030 26880
rect 459646 26868 459652 26880
rect 459704 26868 459710 26920
rect 466822 26868 466828 26920
rect 466880 26908 466886 26920
rect 540974 26908 540980 26920
rect 466880 26880 540980 26908
rect 466880 26868 466886 26880
rect 540974 26868 540980 26880
rect 541032 26868 541038 26920
rect 134058 25576 134064 25628
rect 134116 25616 134122 25628
rect 180886 25616 180892 25628
rect 134116 25588 180892 25616
rect 134116 25576 134122 25588
rect 180886 25576 180892 25588
rect 180944 25576 180950 25628
rect 69014 25508 69020 25560
rect 69072 25548 69078 25560
rect 136634 25548 136640 25560
rect 69072 25520 136640 25548
rect 69072 25508 69078 25520
rect 136634 25508 136640 25520
rect 136692 25508 136698 25560
rect 367094 25508 367100 25560
rect 367152 25548 367158 25560
rect 398834 25548 398840 25560
rect 367152 25520 398840 25548
rect 367152 25508 367158 25520
rect 398834 25508 398840 25520
rect 398892 25508 398898 25560
rect 407206 25508 407212 25560
rect 407264 25548 407270 25560
rect 456886 25548 456892 25560
rect 407264 25520 456892 25548
rect 407264 25508 407270 25520
rect 456886 25508 456892 25520
rect 456944 25508 456950 25560
rect 462314 25508 462320 25560
rect 462372 25548 462378 25560
rect 534074 25548 534080 25560
rect 462372 25520 534080 25548
rect 462372 25508 462378 25520
rect 534074 25508 534080 25520
rect 534132 25508 534138 25560
rect 55214 24080 55220 24132
rect 55272 24120 55278 24132
rect 126974 24120 126980 24132
rect 55272 24092 126980 24120
rect 55272 24080 55278 24092
rect 126974 24080 126980 24092
rect 127032 24080 127038 24132
rect 127066 24080 127072 24132
rect 127124 24120 127130 24132
rect 176746 24120 176752 24132
rect 127124 24092 176752 24120
rect 127124 24080 127130 24092
rect 176746 24080 176752 24092
rect 176804 24080 176810 24132
rect 404446 24080 404452 24132
rect 404504 24120 404510 24132
rect 452746 24120 452752 24132
rect 404504 24092 452752 24120
rect 404504 24080 404510 24092
rect 452746 24080 452752 24092
rect 452804 24080 452810 24132
rect 456978 24080 456984 24132
rect 457036 24120 457042 24132
rect 527174 24120 527180 24132
rect 457036 24092 527180 24120
rect 457036 24080 457042 24092
rect 527174 24080 527180 24092
rect 527232 24080 527238 24132
rect 420914 22788 420920 22840
rect 420972 22828 420978 22840
rect 476206 22828 476212 22840
rect 420972 22800 476212 22828
rect 420972 22788 420978 22800
rect 476206 22788 476212 22800
rect 476264 22788 476270 22840
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 116026 22760 116032 22772
rect 40092 22732 116032 22760
rect 40092 22720 40098 22732
rect 116026 22720 116032 22732
rect 116084 22720 116090 22772
rect 129826 22720 129832 22772
rect 129884 22760 129890 22772
rect 179414 22760 179420 22772
rect 129884 22732 179420 22760
rect 129884 22720 129890 22732
rect 179414 22720 179420 22732
rect 179472 22720 179478 22772
rect 365714 22720 365720 22772
rect 365772 22760 365778 22772
rect 396258 22760 396264 22772
rect 365772 22732 396264 22760
rect 365772 22720 365778 22732
rect 396258 22720 396264 22732
rect 396316 22720 396322 22772
rect 456058 22720 456064 22772
rect 456116 22760 456122 22772
rect 514754 22760 514760 22772
rect 456116 22732 514760 22760
rect 456116 22720 456122 22732
rect 514754 22720 514760 22732
rect 514812 22720 514818 22772
rect 175918 21428 175924 21480
rect 175976 21468 175982 21480
rect 209866 21468 209872 21480
rect 175976 21440 209872 21468
rect 175976 21428 175982 21440
rect 209866 21428 209872 21440
rect 209924 21428 209930 21480
rect 22094 21360 22100 21412
rect 22152 21400 22158 21412
rect 103514 21400 103520 21412
rect 22152 21372 103520 21400
rect 22152 21360 22158 21372
rect 103514 21360 103520 21372
rect 103572 21360 103578 21412
rect 103606 21360 103612 21412
rect 103664 21400 103670 21412
rect 160094 21400 160100 21412
rect 103664 21372 160100 21400
rect 103664 21360 103670 21372
rect 160094 21360 160100 21372
rect 160152 21360 160158 21412
rect 161566 21360 161572 21412
rect 161624 21400 161630 21412
rect 201586 21400 201592 21412
rect 161624 21372 201592 21400
rect 161624 21360 161630 21372
rect 201586 21360 201592 21372
rect 201644 21360 201650 21412
rect 378134 21360 378140 21412
rect 378192 21400 378198 21412
rect 414106 21400 414112 21412
rect 378192 21372 414112 21400
rect 378192 21360 378198 21372
rect 414106 21360 414112 21372
rect 414164 21360 414170 21412
rect 419534 21360 419540 21412
rect 419592 21400 419598 21412
rect 473538 21400 473544 21412
rect 419592 21372 473544 21400
rect 419592 21360 419598 21372
rect 473538 21360 473544 21372
rect 473596 21360 473602 21412
rect 474826 21360 474832 21412
rect 474884 21400 474890 21412
rect 552014 21400 552020 21412
rect 474884 21372 552020 21400
rect 474884 21360 474890 21372
rect 552014 21360 552020 21372
rect 552072 21360 552078 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 511994 20652 512000 20664
rect 3476 20624 512000 20652
rect 3476 20612 3482 20624
rect 511994 20612 512000 20624
rect 512052 20612 512058 20664
rect 577682 20612 577688 20664
rect 577740 20652 577746 20664
rect 579798 20652 579804 20664
rect 577740 20624 579804 20652
rect 577740 20612 577746 20624
rect 579798 20612 579804 20624
rect 579856 20612 579862 20664
rect 157334 18640 157340 18692
rect 157392 18680 157398 18692
rect 197446 18680 197452 18692
rect 157392 18652 197452 18680
rect 157392 18640 157398 18652
rect 197446 18640 197452 18652
rect 197504 18640 197510 18692
rect 372614 18640 372620 18692
rect 372672 18680 372678 18692
rect 407206 18680 407212 18692
rect 372672 18652 407212 18680
rect 372672 18640 372678 18652
rect 407206 18640 407212 18652
rect 407264 18640 407270 18692
rect 100754 18572 100760 18624
rect 100812 18612 100818 18624
rect 158714 18612 158720 18624
rect 100812 18584 158720 18612
rect 100812 18572 100818 18584
rect 158714 18572 158720 18584
rect 158772 18572 158778 18624
rect 392026 18572 392032 18624
rect 392084 18612 392090 18624
rect 434806 18612 434812 18624
rect 392084 18584 434812 18612
rect 392084 18572 392090 18584
rect 434806 18572 434812 18584
rect 434864 18572 434870 18624
rect 451274 18572 451280 18624
rect 451332 18612 451338 18624
rect 518894 18612 518900 18624
rect 451332 18584 518900 18612
rect 451332 18572 451338 18584
rect 518894 18572 518900 18584
rect 518952 18572 518958 18624
rect 399478 17348 399484 17400
rect 399536 17388 399542 17400
rect 441706 17388 441712 17400
rect 399536 17360 441712 17388
rect 399536 17348 399542 17360
rect 441706 17348 441712 17360
rect 441764 17348 441770 17400
rect 162854 17280 162860 17332
rect 162912 17320 162918 17332
rect 201494 17320 201500 17332
rect 162912 17292 201500 17320
rect 162912 17280 162918 17292
rect 201494 17280 201500 17292
rect 201552 17280 201558 17332
rect 57974 17212 57980 17264
rect 58032 17252 58038 17264
rect 128354 17252 128360 17264
rect 58032 17224 128360 17252
rect 58032 17212 58038 17224
rect 128354 17212 128360 17224
rect 128412 17212 128418 17264
rect 143626 17212 143632 17264
rect 143684 17252 143690 17264
rect 187878 17252 187884 17264
rect 143684 17224 187884 17252
rect 143684 17212 143690 17224
rect 187878 17212 187884 17224
rect 187936 17212 187942 17264
rect 383654 17212 383660 17264
rect 383712 17252 383718 17264
rect 423674 17252 423680 17264
rect 383712 17224 423680 17252
rect 383712 17212 383718 17224
rect 423674 17212 423680 17224
rect 423732 17212 423738 17264
rect 441798 17212 441804 17264
rect 441856 17252 441862 17264
rect 505094 17252 505100 17264
rect 441856 17224 505100 17252
rect 441856 17212 441862 17224
rect 505094 17212 505100 17224
rect 505152 17212 505158 17264
rect 158898 15988 158904 16040
rect 158956 16028 158962 16040
rect 198826 16028 198832 16040
rect 158956 16000 198832 16028
rect 158956 15988 158962 16000
rect 198826 15988 198832 16000
rect 198884 15988 198890 16040
rect 139578 15920 139584 15972
rect 139636 15960 139642 15972
rect 185302 15960 185308 15972
rect 139636 15932 185308 15960
rect 139636 15920 139642 15932
rect 185302 15920 185308 15932
rect 185360 15920 185366 15972
rect 427814 15920 427820 15972
rect 427872 15960 427878 15972
rect 484762 15960 484768 15972
rect 427872 15932 484768 15960
rect 427872 15920 427878 15932
rect 484762 15920 484768 15932
rect 484820 15920 484826 15972
rect 51074 15852 51080 15904
rect 51132 15892 51138 15904
rect 122834 15892 122840 15904
rect 51132 15864 122840 15892
rect 51132 15852 51138 15864
rect 122834 15852 122840 15864
rect 122892 15852 122898 15904
rect 123018 15852 123024 15904
rect 123076 15892 123082 15904
rect 173894 15892 173900 15904
rect 123076 15864 173900 15892
rect 123076 15852 123082 15864
rect 173894 15852 173900 15864
rect 173952 15852 173958 15904
rect 329834 15852 329840 15904
rect 329892 15892 329898 15904
rect 345290 15892 345296 15904
rect 329892 15864 345296 15892
rect 329892 15852 329898 15864
rect 345290 15852 345296 15864
rect 345348 15852 345354 15904
rect 353294 15852 353300 15904
rect 353352 15892 353358 15904
rect 378410 15892 378416 15904
rect 353352 15864 378416 15892
rect 353352 15852 353358 15864
rect 378410 15852 378416 15864
rect 378468 15852 378474 15904
rect 389174 15852 389180 15904
rect 389232 15892 389238 15904
rect 430850 15892 430856 15904
rect 389232 15864 430856 15892
rect 389232 15852 389238 15864
rect 430850 15852 430856 15864
rect 430908 15852 430914 15904
rect 459554 15852 459560 15904
rect 459612 15892 459618 15904
rect 531314 15892 531320 15904
rect 459612 15864 531320 15892
rect 459612 15852 459618 15864
rect 531314 15852 531320 15864
rect 531372 15852 531378 15904
rect 386506 14560 386512 14612
rect 386564 14600 386570 14612
rect 426802 14600 426808 14612
rect 386564 14572 426808 14600
rect 386564 14560 386570 14572
rect 426802 14560 426808 14572
rect 426860 14560 426866 14612
rect 422386 14492 422392 14544
rect 422444 14532 422450 14544
rect 478138 14532 478144 14544
rect 422444 14504 478144 14532
rect 422444 14492 422450 14504
rect 478138 14492 478144 14504
rect 478196 14492 478202 14544
rect 69106 14424 69112 14476
rect 69164 14464 69170 14476
rect 135254 14464 135260 14476
rect 69164 14436 135260 14464
rect 69164 14424 69170 14436
rect 135254 14424 135260 14436
rect 135312 14424 135318 14476
rect 135806 14424 135812 14476
rect 135864 14464 135870 14476
rect 183554 14464 183560 14476
rect 135864 14436 183560 14464
rect 135864 14424 135870 14436
rect 183554 14424 183560 14436
rect 183612 14424 183618 14476
rect 183738 14424 183744 14476
rect 183796 14464 183802 14476
rect 216674 14464 216680 14476
rect 183796 14436 216680 14464
rect 183796 14424 183802 14436
rect 216674 14424 216680 14436
rect 216732 14424 216738 14476
rect 345106 14424 345112 14476
rect 345164 14464 345170 14476
rect 367738 14464 367744 14476
rect 345164 14436 367744 14464
rect 345164 14424 345170 14436
rect 367738 14424 367744 14436
rect 367796 14424 367802 14476
rect 394786 14424 394792 14476
rect 394844 14464 394850 14476
rect 439130 14464 439136 14476
rect 394844 14436 439136 14464
rect 394844 14424 394850 14436
rect 439130 14424 439136 14436
rect 439188 14424 439194 14476
rect 476114 14424 476120 14476
rect 476172 14464 476178 14476
rect 554774 14464 554780 14476
rect 476172 14436 554780 14464
rect 476172 14424 476178 14436
rect 554774 14424 554780 14436
rect 554832 14424 554838 14476
rect 351178 13336 351184 13388
rect 351236 13376 351242 13388
rect 371326 13376 371332 13388
rect 351236 13348 371332 13376
rect 351236 13336 351242 13348
rect 371326 13336 371332 13348
rect 371384 13336 371390 13388
rect 371602 13200 371608 13252
rect 371660 13240 371666 13252
rect 406010 13240 406016 13252
rect 371660 13212 406016 13240
rect 371660 13200 371666 13212
rect 406010 13200 406016 13212
rect 406068 13200 406074 13252
rect 150618 13132 150624 13184
rect 150676 13172 150682 13184
rect 193306 13172 193312 13184
rect 150676 13144 193312 13172
rect 150676 13132 150682 13144
rect 193306 13132 193312 13144
rect 193364 13132 193370 13184
rect 387794 13132 387800 13184
rect 387852 13172 387858 13184
rect 428458 13172 428464 13184
rect 387852 13144 428464 13172
rect 387852 13132 387858 13144
rect 428458 13132 428464 13144
rect 428516 13132 428522 13184
rect 132954 13064 132960 13116
rect 133012 13104 133018 13116
rect 180794 13104 180800 13116
rect 133012 13076 180800 13104
rect 133012 13064 133018 13076
rect 180794 13064 180800 13076
rect 180852 13064 180858 13116
rect 205082 13064 205088 13116
rect 205140 13104 205146 13116
rect 230566 13104 230572 13116
rect 205140 13076 230572 13104
rect 205140 13064 205146 13076
rect 230566 13064 230572 13076
rect 230624 13064 230630 13116
rect 360194 13064 360200 13116
rect 360252 13104 360258 13116
rect 389450 13104 389456 13116
rect 360252 13076 389456 13104
rect 360252 13064 360258 13076
rect 389450 13064 389456 13076
rect 389508 13064 389514 13116
rect 403066 13064 403072 13116
rect 403124 13104 403130 13116
rect 449802 13104 449808 13116
rect 403124 13076 449808 13104
rect 403124 13064 403130 13076
rect 449802 13064 449808 13076
rect 449860 13064 449866 13116
rect 470594 13064 470600 13116
rect 470652 13104 470658 13116
rect 547966 13104 547972 13116
rect 470652 13076 547972 13104
rect 470652 13064 470658 13076
rect 547966 13064 547972 13076
rect 548024 13064 548030 13116
rect 345658 12996 345664 13048
rect 345716 13036 345722 13048
rect 353570 13036 353576 13048
rect 345716 13008 353576 13036
rect 345716 12996 345722 13008
rect 353570 12996 353576 13008
rect 353628 12996 353634 13048
rect 338114 11840 338120 11892
rect 338172 11880 338178 11892
rect 357526 11880 357532 11892
rect 338172 11852 357532 11880
rect 338172 11840 338178 11852
rect 357526 11840 357532 11852
rect 357584 11840 357590 11892
rect 137186 11772 137192 11824
rect 137244 11812 137250 11824
rect 183830 11812 183836 11824
rect 137244 11784 183836 11812
rect 137244 11772 137250 11784
rect 183830 11772 183836 11784
rect 183888 11772 183894 11824
rect 342346 11772 342352 11824
rect 342404 11812 342410 11824
rect 364610 11812 364616 11824
rect 342404 11784 364616 11812
rect 342404 11772 342410 11784
rect 364610 11772 364616 11784
rect 364668 11772 364674 11824
rect 367278 11772 367284 11824
rect 367336 11812 367342 11824
rect 399018 11812 399024 11824
rect 367336 11784 399024 11812
rect 367336 11772 367342 11784
rect 399018 11772 399024 11784
rect 399076 11772 399082 11824
rect 24210 11704 24216 11756
rect 24268 11744 24274 11756
rect 104158 11744 104164 11756
rect 24268 11716 104164 11744
rect 24268 11704 24274 11716
rect 104158 11704 104164 11716
rect 104216 11704 104222 11756
rect 128906 11704 128912 11756
rect 128964 11744 128970 11756
rect 178126 11744 178132 11756
rect 128964 11716 178132 11744
rect 128964 11704 128970 11716
rect 178126 11704 178132 11716
rect 178184 11704 178190 11756
rect 186130 11704 186136 11756
rect 186188 11744 186194 11756
rect 218054 11744 218060 11756
rect 186188 11716 218060 11744
rect 186188 11704 186194 11716
rect 218054 11704 218060 11716
rect 218112 11704 218118 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 259454 11704 259460 11756
rect 259512 11744 259518 11756
rect 260650 11744 260656 11756
rect 259512 11716 260656 11744
rect 259512 11704 259518 11716
rect 260650 11704 260656 11716
rect 260708 11704 260714 11756
rect 356698 11704 356704 11756
rect 356756 11744 356762 11756
rect 382366 11744 382372 11756
rect 356756 11716 382372 11744
rect 356756 11704 356762 11716
rect 382366 11704 382372 11716
rect 382424 11704 382430 11756
rect 391934 11704 391940 11756
rect 391992 11744 391998 11756
rect 433978 11744 433984 11756
rect 391992 11716 433984 11744
rect 391992 11704 391998 11716
rect 433978 11704 433984 11716
rect 434036 11704 434042 11756
rect 438946 11704 438952 11756
rect 439004 11744 439010 11756
rect 501322 11744 501328 11756
rect 439004 11716 501328 11744
rect 439004 11704 439010 11716
rect 501322 11704 501328 11716
rect 501380 11704 501386 11756
rect 363598 10412 363604 10464
rect 363656 10452 363662 10464
rect 391106 10452 391112 10464
rect 363656 10424 391112 10452
rect 363656 10412 363662 10424
rect 391106 10412 391112 10424
rect 391164 10412 391170 10464
rect 111610 10344 111616 10396
rect 111668 10384 111674 10396
rect 165706 10384 165712 10396
rect 111668 10356 165712 10384
rect 111668 10344 111674 10356
rect 165706 10344 165712 10356
rect 165764 10344 165770 10396
rect 178678 10344 178684 10396
rect 178736 10384 178742 10396
rect 211246 10384 211252 10396
rect 178736 10356 211252 10384
rect 178736 10344 178742 10356
rect 211246 10344 211252 10356
rect 211304 10344 211310 10396
rect 332686 10344 332692 10396
rect 332744 10384 332750 10396
rect 349154 10384 349160 10396
rect 332744 10356 349160 10384
rect 332744 10344 332750 10356
rect 349154 10344 349160 10356
rect 349212 10344 349218 10396
rect 364426 10344 364432 10396
rect 364484 10384 364490 10396
rect 395338 10384 395344 10396
rect 364484 10356 395344 10384
rect 364484 10344 364490 10356
rect 395338 10344 395344 10356
rect 395396 10344 395402 10396
rect 429194 10344 429200 10396
rect 429252 10384 429258 10396
rect 487154 10384 487160 10396
rect 429252 10356 487160 10384
rect 429252 10344 429258 10356
rect 487154 10344 487160 10356
rect 487212 10344 487218 10396
rect 65058 10276 65064 10328
rect 65116 10316 65122 10328
rect 133874 10316 133880 10328
rect 65116 10288 133880 10316
rect 65116 10276 65122 10288
rect 133874 10276 133880 10288
rect 133932 10276 133938 10328
rect 164418 10276 164424 10328
rect 164476 10316 164482 10328
rect 202874 10316 202880 10328
rect 164476 10288 202880 10316
rect 164476 10276 164482 10288
rect 202874 10276 202880 10288
rect 202932 10276 202938 10328
rect 342254 10276 342260 10328
rect 342312 10316 342318 10328
rect 363506 10316 363512 10328
rect 342312 10288 363512 10316
rect 342312 10276 342318 10288
rect 363506 10276 363512 10288
rect 363564 10276 363570 10328
rect 378226 10276 378232 10328
rect 378284 10316 378290 10328
rect 415486 10316 415492 10328
rect 378284 10288 415492 10316
rect 378284 10276 378290 10288
rect 415486 10276 415492 10288
rect 415544 10276 415550 10328
rect 473446 10276 473452 10328
rect 473504 10316 473510 10328
rect 551002 10316 551008 10328
rect 473504 10288 551008 10316
rect 473504 10276 473510 10288
rect 551002 10276 551008 10288
rect 551060 10276 551066 10328
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 161290 9052 161296 9104
rect 161348 9092 161354 9104
rect 200206 9092 200212 9104
rect 161348 9064 200212 9092
rect 161348 9052 161354 9064
rect 200206 9052 200212 9064
rect 200264 9052 200270 9104
rect 358814 9052 358820 9104
rect 358872 9092 358878 9104
rect 388254 9092 388260 9104
rect 358872 9064 388260 9092
rect 358872 9052 358878 9064
rect 388254 9052 388260 9064
rect 388312 9052 388318 9104
rect 109310 8984 109316 9036
rect 109368 9024 109374 9036
rect 164326 9024 164332 9036
rect 109368 8996 164332 9024
rect 109368 8984 109374 8996
rect 164326 8984 164332 8996
rect 164384 8984 164390 9036
rect 169570 8984 169576 9036
rect 169628 9024 169634 9036
rect 206002 9024 206008 9036
rect 169628 8996 206008 9024
rect 169628 8984 169634 8996
rect 206002 8984 206008 8996
rect 206060 8984 206066 9036
rect 328454 8984 328460 9036
rect 328512 9024 328518 9036
rect 343358 9024 343364 9036
rect 328512 8996 343364 9024
rect 328512 8984 328518 8996
rect 343358 8984 343364 8996
rect 343416 8984 343422 9036
rect 382274 8984 382280 9036
rect 382332 9024 382338 9036
rect 420178 9024 420184 9036
rect 382332 8996 420184 9024
rect 382332 8984 382338 8996
rect 420178 8984 420184 8996
rect 420236 8984 420242 9036
rect 426434 8984 426440 9036
rect 426492 9024 426498 9036
rect 484026 9024 484032 9036
rect 426492 8996 484032 9024
rect 426492 8984 426498 8996
rect 484026 8984 484032 8996
rect 484084 8984 484090 9036
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 110414 8956 110420 8968
rect 33652 8928 110420 8956
rect 33652 8916 33658 8928
rect 110414 8916 110420 8928
rect 110472 8916 110478 8968
rect 128170 8916 128176 8968
rect 128228 8956 128234 8968
rect 176654 8956 176660 8968
rect 128228 8928 176660 8956
rect 128228 8916 128234 8928
rect 176654 8916 176660 8928
rect 176712 8916 176718 8968
rect 336826 8916 336832 8968
rect 336884 8956 336890 8968
rect 356330 8956 356336 8968
rect 336884 8928 356336 8956
rect 336884 8916 336890 8928
rect 356330 8916 356336 8928
rect 356388 8916 356394 8968
rect 359458 8916 359464 8968
rect 359516 8956 359522 8968
rect 384758 8956 384764 8968
rect 359516 8928 384764 8956
rect 359516 8916 359522 8928
rect 384758 8916 384764 8928
rect 384816 8916 384822 8968
rect 385126 8916 385132 8968
rect 385184 8956 385190 8968
rect 424962 8956 424968 8968
rect 385184 8928 424968 8956
rect 385184 8916 385190 8928
rect 424962 8916 424968 8928
rect 425020 8916 425026 8968
rect 454034 8916 454040 8968
rect 454092 8956 454098 8968
rect 523034 8956 523040 8968
rect 454092 8928 523040 8956
rect 454092 8916 454098 8928
rect 523034 8916 523040 8928
rect 523092 8916 523098 8968
rect 351914 7760 351920 7812
rect 351972 7800 351978 7812
rect 377674 7800 377680 7812
rect 351972 7772 377680 7800
rect 351972 7760 351978 7772
rect 377674 7760 377680 7772
rect 377732 7760 377738 7812
rect 321646 7692 321652 7744
rect 321704 7732 321710 7744
rect 335078 7732 335084 7744
rect 321704 7704 335084 7732
rect 321704 7692 321710 7704
rect 335078 7692 335084 7704
rect 335136 7692 335142 7744
rect 354674 7692 354680 7744
rect 354732 7732 354738 7744
rect 381170 7732 381176 7744
rect 354732 7704 381176 7732
rect 354732 7692 354738 7704
rect 381170 7692 381176 7704
rect 381228 7692 381234 7744
rect 125870 7624 125876 7676
rect 125928 7664 125934 7676
rect 175366 7664 175372 7676
rect 125928 7636 175372 7664
rect 125928 7624 125934 7636
rect 175366 7624 175372 7636
rect 175424 7624 175430 7676
rect 203886 7624 203892 7676
rect 203944 7664 203950 7676
rect 230474 7664 230480 7676
rect 203944 7636 230480 7664
rect 203944 7624 203950 7636
rect 230474 7624 230480 7636
rect 230532 7624 230538 7676
rect 331858 7624 331864 7676
rect 331916 7664 331922 7676
rect 346946 7664 346952 7676
rect 331916 7636 346952 7664
rect 331916 7624 331922 7636
rect 346946 7624 346952 7636
rect 347004 7624 347010 7676
rect 379514 7624 379520 7676
rect 379572 7664 379578 7676
rect 416682 7664 416688 7676
rect 379572 7636 416688 7664
rect 379572 7624 379578 7636
rect 416682 7624 416688 7636
rect 416740 7624 416746 7676
rect 448606 7624 448612 7676
rect 448664 7664 448670 7676
rect 515950 7664 515956 7676
rect 448664 7636 515956 7664
rect 448664 7624 448670 7636
rect 515950 7624 515956 7636
rect 516008 7624 516014 7676
rect 7650 7556 7656 7608
rect 7708 7596 7714 7608
rect 92566 7596 92572 7608
rect 7708 7568 92572 7596
rect 7708 7556 7714 7568
rect 92566 7556 92572 7568
rect 92624 7556 92630 7608
rect 105722 7556 105728 7608
rect 105780 7596 105786 7608
rect 161474 7596 161480 7608
rect 105780 7568 161480 7596
rect 105780 7556 105786 7568
rect 161474 7556 161480 7568
rect 161532 7556 161538 7608
rect 168374 7556 168380 7608
rect 168432 7596 168438 7608
rect 205726 7596 205732 7608
rect 168432 7568 205732 7596
rect 168432 7556 168438 7568
rect 205726 7556 205732 7568
rect 205784 7556 205790 7608
rect 334342 7556 334348 7608
rect 334400 7596 334406 7608
rect 352834 7596 352840 7608
rect 334400 7568 352840 7596
rect 334400 7556 334406 7568
rect 352834 7556 352840 7568
rect 352892 7556 352898 7608
rect 376846 7556 376852 7608
rect 376904 7596 376910 7608
rect 413094 7596 413100 7608
rect 376904 7568 413100 7596
rect 376904 7556 376910 7568
rect 413094 7556 413100 7568
rect 413152 7556 413158 7608
rect 423858 7556 423864 7608
rect 423916 7596 423922 7608
rect 480530 7596 480536 7608
rect 423916 7568 480536 7596
rect 423916 7556 423922 7568
rect 480530 7556 480536 7568
rect 480588 7556 480594 7608
rect 485866 7556 485872 7608
rect 485924 7596 485930 7608
rect 569126 7596 569132 7608
rect 485924 7568 569132 7596
rect 485924 7556 485930 7568
rect 569126 7556 569132 7568
rect 569184 7556 569190 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 511074 6848 511080 6860
rect 3476 6820 511080 6848
rect 3476 6808 3482 6820
rect 511074 6808 511080 6820
rect 511132 6808 511138 6860
rect 577498 6740 577504 6792
rect 577556 6780 577562 6792
rect 579706 6780 579712 6792
rect 577556 6752 579712 6780
rect 577556 6740 577562 6752
rect 579706 6740 579712 6752
rect 579764 6740 579770 6792
rect 77386 6604 77392 6656
rect 77444 6644 77450 6656
rect 142154 6644 142160 6656
rect 77444 6616 142160 6644
rect 77444 6604 77450 6616
rect 142154 6604 142160 6616
rect 142212 6604 142218 6656
rect 434714 6604 434720 6656
rect 434772 6644 434778 6656
rect 495894 6644 495900 6656
rect 434772 6616 495900 6644
rect 434772 6604 434778 6616
rect 495894 6604 495900 6616
rect 495952 6604 495958 6656
rect 66714 6536 66720 6588
rect 66772 6576 66778 6588
rect 134150 6576 134156 6588
rect 66772 6548 134156 6576
rect 66772 6536 66778 6548
rect 134150 6536 134156 6548
rect 134208 6536 134214 6588
rect 437474 6536 437480 6588
rect 437532 6576 437538 6588
rect 499390 6576 499396 6588
rect 437532 6548 499396 6576
rect 437532 6536 437538 6548
rect 499390 6536 499396 6548
rect 499448 6536 499454 6588
rect 63218 6468 63224 6520
rect 63276 6508 63282 6520
rect 131114 6508 131120 6520
rect 63276 6480 131120 6508
rect 63276 6468 63282 6480
rect 131114 6468 131120 6480
rect 131172 6468 131178 6520
rect 440234 6468 440240 6520
rect 440292 6508 440298 6520
rect 502978 6508 502984 6520
rect 440292 6480 502984 6508
rect 440292 6468 440298 6480
rect 502978 6468 502984 6480
rect 503036 6468 503042 6520
rect 59630 6400 59636 6452
rect 59688 6440 59694 6452
rect 129734 6440 129740 6452
rect 59688 6412 129740 6440
rect 59688 6400 59694 6412
rect 129734 6400 129740 6412
rect 129792 6400 129798 6452
rect 346486 6400 346492 6452
rect 346544 6440 346550 6452
rect 370590 6440 370596 6452
rect 346544 6412 370596 6440
rect 346544 6400 346550 6412
rect 370590 6400 370596 6412
rect 370648 6400 370654 6452
rect 444466 6400 444472 6452
rect 444524 6440 444530 6452
rect 510062 6440 510068 6452
rect 444524 6412 510068 6440
rect 444524 6400 444530 6412
rect 510062 6400 510068 6412
rect 510120 6400 510126 6452
rect 52546 6332 52552 6384
rect 52604 6372 52610 6384
rect 124306 6372 124312 6384
rect 52604 6344 124312 6372
rect 52604 6332 52610 6344
rect 124306 6332 124312 6344
rect 124364 6332 124370 6384
rect 441614 6332 441620 6384
rect 441672 6372 441678 6384
rect 506474 6372 506480 6384
rect 441672 6344 506480 6372
rect 441672 6332 441678 6344
rect 506474 6332 506480 6344
rect 506532 6332 506538 6384
rect 48958 6264 48964 6316
rect 49016 6304 49022 6316
rect 121730 6304 121736 6316
rect 49016 6276 121736 6304
rect 49016 6264 49022 6276
rect 121730 6264 121736 6276
rect 121788 6264 121794 6316
rect 138842 6264 138848 6316
rect 138900 6304 138906 6316
rect 185026 6304 185032 6316
rect 138900 6276 185032 6304
rect 138900 6264 138906 6276
rect 185026 6264 185032 6276
rect 185084 6264 185090 6316
rect 370038 6264 370044 6316
rect 370096 6304 370102 6316
rect 402514 6304 402520 6316
rect 370096 6276 402520 6304
rect 370096 6264 370102 6276
rect 402514 6264 402520 6276
rect 402572 6264 402578 6316
rect 449894 6264 449900 6316
rect 449952 6304 449958 6316
rect 517146 6304 517152 6316
rect 449952 6276 517152 6304
rect 449952 6264 449958 6276
rect 517146 6264 517152 6276
rect 517204 6264 517210 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 93946 6236 93952 6248
rect 8812 6208 93952 6236
rect 8812 6196 8818 6208
rect 93946 6196 93952 6208
rect 94004 6196 94010 6248
rect 131758 6196 131764 6248
rect 131816 6236 131822 6248
rect 179598 6236 179604 6248
rect 131816 6208 179604 6236
rect 131816 6196 131822 6208
rect 179598 6196 179604 6208
rect 179656 6196 179662 6248
rect 213362 6196 213368 6248
rect 213420 6236 213426 6248
rect 237374 6236 237380 6248
rect 213420 6208 237380 6236
rect 213420 6196 213426 6208
rect 237374 6196 237380 6208
rect 237432 6196 237438 6248
rect 374178 6196 374184 6248
rect 374236 6236 374242 6248
rect 409598 6236 409604 6248
rect 374236 6208 409604 6236
rect 374236 6196 374242 6208
rect 409598 6196 409604 6208
rect 409656 6196 409662 6248
rect 447134 6196 447140 6248
rect 447192 6236 447198 6248
rect 513558 6236 513564 6248
rect 447192 6208 513564 6236
rect 447192 6196 447198 6208
rect 513558 6196 513564 6208
rect 513616 6196 513622 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 89714 6168 89720 6180
rect 4120 6140 89720 6168
rect 4120 6128 4126 6140
rect 89714 6128 89720 6140
rect 89772 6128 89778 6180
rect 118786 6128 118792 6180
rect 118844 6168 118850 6180
rect 171226 6168 171232 6180
rect 118844 6140 171232 6168
rect 118844 6128 118850 6140
rect 171226 6128 171232 6140
rect 171284 6128 171290 6180
rect 182542 6128 182548 6180
rect 182600 6168 182606 6180
rect 215294 6168 215300 6180
rect 182600 6140 215300 6168
rect 182600 6128 182606 6140
rect 215294 6128 215300 6140
rect 215352 6128 215358 6180
rect 327074 6128 327080 6180
rect 327132 6168 327138 6180
rect 342162 6168 342168 6180
rect 327132 6140 342168 6168
rect 327132 6128 327138 6140
rect 342162 6128 342168 6140
rect 342220 6128 342226 6180
rect 349246 6128 349252 6180
rect 349304 6168 349310 6180
rect 374086 6168 374092 6180
rect 349304 6140 374092 6168
rect 349304 6128 349310 6140
rect 374086 6128 374092 6140
rect 374144 6128 374150 6180
rect 388162 6128 388168 6180
rect 388220 6168 388226 6180
rect 429654 6168 429660 6180
rect 388220 6140 429660 6168
rect 388220 6128 388226 6140
rect 429654 6128 429660 6140
rect 429712 6128 429718 6180
rect 452654 6128 452660 6180
rect 452712 6168 452718 6180
rect 520734 6168 520740 6180
rect 452712 6140 520740 6168
rect 452712 6128 452718 6140
rect 520734 6128 520740 6140
rect 520792 6128 520798 6180
rect 336090 5516 336096 5568
rect 336148 5556 336154 5568
rect 339862 5556 339868 5568
rect 336148 5528 339868 5556
rect 336148 5516 336154 5528
rect 339862 5516 339868 5528
rect 339920 5516 339926 5568
rect 93946 5380 93952 5432
rect 94004 5420 94010 5432
rect 153194 5420 153200 5432
rect 94004 5392 153200 5420
rect 94004 5380 94010 5392
rect 153194 5380 153200 5392
rect 153252 5380 153258 5432
rect 90358 5312 90364 5364
rect 90416 5352 90422 5364
rect 150710 5352 150716 5364
rect 90416 5324 150716 5352
rect 90416 5312 90422 5324
rect 150710 5312 150716 5324
rect 150768 5312 150774 5364
rect 394694 5312 394700 5364
rect 394752 5352 394758 5364
rect 437934 5352 437940 5364
rect 394752 5324 437940 5352
rect 394752 5312 394758 5324
rect 437934 5312 437940 5324
rect 437992 5312 437998 5364
rect 86862 5244 86868 5296
rect 86920 5284 86926 5296
rect 147674 5284 147680 5296
rect 86920 5256 147680 5284
rect 86920 5244 86926 5256
rect 147674 5244 147680 5256
rect 147732 5244 147738 5296
rect 396166 5244 396172 5296
rect 396224 5284 396230 5296
rect 441522 5284 441528 5296
rect 396224 5256 441528 5284
rect 396224 5244 396230 5256
rect 441522 5244 441528 5256
rect 441580 5244 441586 5296
rect 456794 5244 456800 5296
rect 456852 5284 456858 5296
rect 526622 5284 526628 5296
rect 456852 5256 526628 5284
rect 456852 5244 456858 5256
rect 526622 5244 526628 5256
rect 526680 5244 526686 5296
rect 83274 5176 83280 5228
rect 83332 5216 83338 5228
rect 146294 5216 146300 5228
rect 83332 5188 146300 5216
rect 83332 5176 83338 5188
rect 146294 5176 146300 5188
rect 146352 5176 146358 5228
rect 398926 5176 398932 5228
rect 398984 5216 398990 5228
rect 445018 5216 445024 5228
rect 398984 5188 445024 5216
rect 398984 5176 398990 5188
rect 445018 5176 445024 5188
rect 445076 5176 445082 5228
rect 461026 5176 461032 5228
rect 461084 5216 461090 5228
rect 533706 5216 533712 5228
rect 461084 5188 533712 5216
rect 461084 5176 461090 5188
rect 533706 5176 533712 5188
rect 533764 5176 533770 5228
rect 79686 5108 79692 5160
rect 79744 5148 79750 5160
rect 143626 5148 143632 5160
rect 79744 5120 143632 5148
rect 79744 5108 79750 5120
rect 143626 5108 143632 5120
rect 143684 5108 143690 5160
rect 404354 5108 404360 5160
rect 404412 5148 404418 5160
rect 452102 5148 452108 5160
rect 404412 5120 452108 5148
rect 404412 5108 404418 5120
rect 452102 5108 452108 5120
rect 452160 5108 452166 5160
rect 458174 5108 458180 5160
rect 458232 5148 458238 5160
rect 530118 5148 530124 5160
rect 458232 5120 530124 5148
rect 458232 5108 458238 5120
rect 530118 5108 530124 5120
rect 530176 5108 530182 5160
rect 76190 5040 76196 5092
rect 76248 5080 76254 5092
rect 140774 5080 140780 5092
rect 76248 5052 140780 5080
rect 76248 5040 76254 5052
rect 140774 5040 140780 5052
rect 140832 5040 140838 5092
rect 407114 5040 407120 5092
rect 407172 5080 407178 5092
rect 455690 5080 455696 5092
rect 407172 5052 455696 5080
rect 407172 5040 407178 5052
rect 455690 5040 455696 5052
rect 455748 5040 455754 5092
rect 466454 5040 466460 5092
rect 466512 5080 466518 5092
rect 540790 5080 540796 5092
rect 466512 5052 540796 5080
rect 466512 5040 466518 5052
rect 540790 5040 540796 5052
rect 540848 5040 540854 5092
rect 72602 4972 72608 5024
rect 72660 5012 72666 5024
rect 138198 5012 138204 5024
rect 72660 4984 138204 5012
rect 72660 4972 72666 4984
rect 138198 4972 138204 4984
rect 138256 4972 138262 5024
rect 154206 4972 154212 5024
rect 154264 5012 154270 5024
rect 195974 5012 195980 5024
rect 154264 4984 195980 5012
rect 154264 4972 154270 4984
rect 195974 4972 195980 4984
rect 196032 4972 196038 5024
rect 408862 4972 408868 5024
rect 408920 5012 408926 5024
rect 459186 5012 459192 5024
rect 408920 4984 459192 5012
rect 408920 4972 408926 4984
rect 459186 4972 459192 4984
rect 459244 4972 459250 5024
rect 463694 4972 463700 5024
rect 463752 5012 463758 5024
rect 537202 5012 537208 5024
rect 463752 4984 537208 5012
rect 463752 4972 463758 4984
rect 537202 4972 537208 4984
rect 537260 4972 537266 5024
rect 21818 4904 21824 4956
rect 21876 4944 21882 4956
rect 102502 4944 102508 4956
rect 21876 4916 102508 4944
rect 21876 4904 21882 4916
rect 102502 4904 102508 4916
rect 102560 4904 102566 4956
rect 144730 4904 144736 4956
rect 144788 4944 144794 4956
rect 189074 4944 189080 4956
rect 144788 4916 189080 4944
rect 144788 4904 144794 4916
rect 189074 4904 189080 4916
rect 189132 4904 189138 4956
rect 314654 4904 314660 4956
rect 314712 4944 314718 4956
rect 324314 4944 324320 4956
rect 314712 4916 324320 4944
rect 314712 4904 314718 4916
rect 324314 4904 324320 4916
rect 324372 4904 324378 4956
rect 349798 4904 349804 4956
rect 349856 4944 349862 4956
rect 367002 4944 367008 4956
rect 349856 4916 367008 4944
rect 349856 4904 349862 4916
rect 367002 4904 367008 4916
rect 367060 4904 367066 4956
rect 411346 4904 411352 4956
rect 411404 4944 411410 4956
rect 462774 4944 462780 4956
rect 411404 4916 462780 4944
rect 411404 4904 411410 4916
rect 462774 4904 462780 4916
rect 462832 4904 462838 4956
rect 469214 4904 469220 4956
rect 469272 4944 469278 4956
rect 544378 4944 544384 4956
rect 469272 4916 544384 4944
rect 469272 4904 469278 4916
rect 544378 4904 544384 4916
rect 544436 4904 544442 4956
rect 17034 4836 17040 4888
rect 17092 4876 17098 4888
rect 99374 4876 99380 4888
rect 17092 4848 99380 4876
rect 17092 4836 17098 4848
rect 99374 4836 99380 4848
rect 99432 4836 99438 4888
rect 141234 4836 141240 4888
rect 141292 4876 141298 4888
rect 186314 4876 186320 4888
rect 141292 4848 186320 4876
rect 141292 4836 141298 4848
rect 186314 4836 186320 4848
rect 186372 4836 186378 4888
rect 241698 4836 241704 4888
rect 241756 4876 241762 4888
rect 256786 4876 256792 4888
rect 241756 4848 256792 4876
rect 241756 4836 241762 4848
rect 256786 4836 256792 4848
rect 256844 4836 256850 4888
rect 332594 4836 332600 4888
rect 332652 4876 332658 4888
rect 349246 4876 349252 4888
rect 332652 4848 349252 4876
rect 332652 4836 332658 4848
rect 349246 4836 349252 4848
rect 349304 4836 349310 4888
rect 355318 4836 355324 4888
rect 355376 4876 355382 4888
rect 375282 4876 375288 4888
rect 355376 4848 375288 4876
rect 355376 4836 355382 4848
rect 375282 4836 375288 4848
rect 375340 4836 375346 4888
rect 414014 4836 414020 4888
rect 414072 4876 414078 4888
rect 466270 4876 466276 4888
rect 414072 4848 466276 4876
rect 414072 4836 414078 4848
rect 466270 4836 466276 4848
rect 466328 4836 466334 4888
rect 491294 4836 491300 4888
rect 491352 4876 491358 4888
rect 576302 4876 576308 4888
rect 491352 4848 576308 4876
rect 491352 4836 491358 4848
rect 576302 4836 576308 4848
rect 576360 4836 576366 4888
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 96614 4808 96620 4820
rect 12400 4780 96620 4808
rect 12400 4768 12406 4780
rect 96614 4768 96620 4780
rect 96672 4768 96678 4820
rect 97442 4768 97448 4820
rect 97500 4808 97506 4820
rect 155954 4808 155960 4820
rect 97500 4780 155960 4808
rect 97500 4768 97506 4780
rect 155954 4768 155960 4780
rect 156012 4768 156018 4820
rect 194410 4768 194416 4820
rect 194468 4808 194474 4820
rect 223574 4808 223580 4820
rect 194468 4780 223580 4808
rect 194468 4768 194474 4780
rect 223574 4768 223580 4780
rect 223632 4768 223638 4820
rect 235810 4768 235816 4820
rect 235868 4808 235874 4820
rect 252554 4808 252560 4820
rect 235868 4780 252560 4808
rect 235868 4768 235874 4780
rect 252554 4768 252560 4780
rect 252612 4768 252618 4820
rect 253474 4768 253480 4820
rect 253532 4808 253538 4820
rect 265066 4808 265072 4820
rect 253532 4780 265072 4808
rect 253532 4768 253538 4780
rect 265066 4768 265072 4780
rect 265124 4768 265130 4820
rect 324406 4768 324412 4820
rect 324464 4808 324470 4820
rect 338666 4808 338672 4820
rect 324464 4780 338672 4808
rect 324464 4768 324470 4780
rect 338666 4768 338672 4780
rect 338724 4768 338730 4820
rect 339586 4768 339592 4820
rect 339644 4808 339650 4820
rect 359918 4808 359924 4820
rect 339644 4780 359924 4808
rect 339644 4768 339650 4780
rect 359918 4768 359924 4780
rect 359976 4768 359982 4820
rect 362954 4768 362960 4820
rect 363012 4808 363018 4820
rect 393038 4808 393044 4820
rect 363012 4780 393044 4808
rect 363012 4768 363018 4780
rect 393038 4768 393044 4780
rect 393096 4768 393102 4820
rect 416774 4768 416780 4820
rect 416832 4808 416838 4820
rect 469858 4808 469864 4820
rect 416832 4780 469864 4808
rect 416832 4768 416838 4780
rect 469858 4768 469864 4780
rect 469916 4768 469922 4820
rect 488534 4768 488540 4820
rect 488592 4808 488598 4820
rect 572714 4808 572720 4820
rect 488592 4780 572720 4808
rect 488592 4768 488598 4780
rect 572714 4768 572720 4780
rect 572772 4768 572778 4820
rect 323578 4360 323584 4412
rect 323636 4400 323642 4412
rect 327994 4400 328000 4412
rect 323636 4372 328000 4400
rect 323636 4360 323642 4372
rect 327994 4360 328000 4372
rect 328052 4360 328058 4412
rect 327718 4156 327724 4208
rect 327776 4196 327782 4208
rect 331582 4196 331588 4208
rect 327776 4168 331588 4196
rect 327776 4156 327782 4168
rect 331582 4156 331588 4168
rect 331640 4156 331646 4208
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 7558 4128 7564 4140
rect 1728 4100 7564 4128
rect 1728 4088 1734 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 17218 4128 17224 4140
rect 13596 4100 17224 4128
rect 13596 4088 13602 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 180242 4088 180248 4140
rect 180300 4128 180306 4140
rect 182818 4128 182824 4140
rect 180300 4100 182824 4128
rect 180300 4088 180306 4100
rect 182818 4088 182824 4100
rect 182876 4088 182882 4140
rect 262950 4088 262956 4140
rect 263008 4128 263014 4140
rect 269758 4128 269764 4140
rect 263008 4100 269764 4128
rect 263008 4088 263014 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 284294 4088 284300 4140
rect 284352 4128 284358 4140
rect 287146 4128 287152 4140
rect 284352 4100 287152 4128
rect 284352 4088 284358 4100
rect 287146 4088 287152 4100
rect 287204 4088 287210 4140
rect 302326 4088 302332 4140
rect 302384 4128 302390 4140
rect 303522 4128 303528 4140
rect 302384 4100 303528 4128
rect 302384 4088 302390 4100
rect 303522 4088 303528 4100
rect 303580 4088 303586 4140
rect 436738 4088 436744 4140
rect 436796 4128 436802 4140
rect 443822 4128 443828 4140
rect 436796 4100 443828 4128
rect 436796 4088 436802 4100
rect 443822 4088 443828 4100
rect 443880 4088 443886 4140
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 28258 4060 28264 4072
rect 20680 4032 28264 4060
rect 20680 4020 20686 4032
rect 28258 4020 28264 4032
rect 28316 4020 28322 4072
rect 208578 4020 208584 4072
rect 208636 4060 208642 4072
rect 221458 4060 221464 4072
rect 208636 4032 221464 4060
rect 208636 4020 208642 4032
rect 221458 4020 221464 4032
rect 221516 4020 221522 4072
rect 201494 3952 201500 4004
rect 201552 3992 201558 4004
rect 217318 3992 217324 4004
rect 201552 3964 217324 3992
rect 201552 3952 201558 3964
rect 217318 3952 217324 3964
rect 217376 3952 217382 4004
rect 398098 3952 398104 4004
rect 398156 3992 398162 4004
rect 408402 3992 408408 4004
rect 398156 3964 408408 3992
rect 398156 3952 398162 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 114002 3884 114008 3936
rect 114060 3924 114066 3936
rect 156598 3924 156604 3936
rect 114060 3896 156604 3924
rect 114060 3884 114066 3896
rect 156598 3884 156604 3896
rect 156656 3884 156662 3936
rect 216858 3884 216864 3936
rect 216916 3924 216922 3936
rect 235258 3924 235264 3936
rect 216916 3896 235264 3924
rect 216916 3884 216922 3896
rect 235258 3884 235264 3896
rect 235316 3884 235322 3936
rect 305638 3884 305644 3936
rect 305696 3924 305702 3936
rect 309042 3924 309048 3936
rect 305696 3896 309048 3924
rect 305696 3884 305702 3896
rect 309042 3884 309048 3896
rect 309100 3884 309106 3936
rect 313918 3884 313924 3936
rect 313976 3924 313982 3936
rect 320910 3924 320916 3936
rect 313976 3896 320916 3924
rect 313976 3884 313982 3896
rect 320910 3884 320916 3896
rect 320968 3884 320974 3936
rect 321554 3884 321560 3936
rect 321612 3924 321618 3936
rect 333882 3924 333888 3936
rect 321612 3896 333888 3924
rect 321612 3884 321618 3896
rect 333882 3884 333888 3896
rect 333940 3884 333946 3936
rect 335998 3884 336004 3936
rect 336056 3924 336062 3936
rect 351638 3924 351644 3936
rect 336056 3896 351644 3924
rect 336056 3884 336062 3896
rect 351638 3884 351644 3896
rect 351696 3884 351702 3936
rect 380894 3884 380900 3936
rect 380952 3924 380958 3936
rect 418982 3924 418988 3936
rect 380952 3896 418988 3924
rect 380952 3884 380958 3896
rect 418982 3884 418988 3896
rect 419040 3884 419046 3936
rect 542998 3884 543004 3936
rect 543056 3924 543062 3936
rect 557350 3924 557356 3936
rect 543056 3896 557356 3924
rect 543056 3884 543062 3896
rect 557350 3884 557356 3896
rect 557408 3884 557414 3936
rect 89162 3816 89168 3868
rect 89220 3856 89226 3868
rect 140038 3856 140044 3868
rect 89220 3828 140044 3856
rect 89220 3816 89226 3828
rect 140038 3816 140044 3828
rect 140096 3816 140102 3868
rect 215662 3816 215668 3868
rect 215720 3856 215726 3868
rect 233878 3856 233884 3868
rect 215720 3828 233884 3856
rect 215720 3816 215726 3828
rect 233878 3816 233884 3828
rect 233936 3816 233942 3868
rect 276014 3816 276020 3868
rect 276072 3856 276078 3868
rect 278038 3856 278044 3868
rect 276072 3828 278044 3856
rect 276072 3816 276078 3828
rect 278038 3816 278044 3828
rect 278096 3816 278102 3868
rect 316126 3816 316132 3868
rect 316184 3856 316190 3868
rect 326798 3856 326804 3868
rect 316184 3828 326804 3856
rect 316184 3816 316190 3828
rect 326798 3816 326804 3828
rect 326856 3816 326862 3868
rect 328546 3816 328552 3868
rect 328604 3856 328610 3868
rect 344554 3856 344560 3868
rect 328604 3828 344560 3856
rect 328604 3816 328610 3828
rect 344554 3816 344560 3828
rect 344612 3816 344618 3868
rect 386414 3816 386420 3868
rect 386472 3856 386478 3868
rect 426158 3856 426164 3868
rect 386472 3828 426164 3856
rect 386472 3816 386478 3828
rect 426158 3816 426164 3828
rect 426216 3816 426222 3868
rect 440878 3816 440884 3868
rect 440936 3856 440942 3868
rect 450906 3856 450912 3868
rect 440936 3828 450912 3856
rect 440936 3816 440942 3828
rect 450906 3816 450912 3828
rect 450964 3816 450970 3868
rect 545758 3816 545764 3868
rect 545816 3856 545822 3868
rect 564434 3856 564440 3868
rect 545816 3828 564440 3856
rect 545816 3816 545822 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 50338 3788 50344 3800
rect 43128 3760 50344 3788
rect 43128 3748 43134 3760
rect 50338 3748 50344 3760
rect 50396 3748 50402 3800
rect 82078 3748 82084 3800
rect 82136 3788 82142 3800
rect 135898 3788 135904 3800
rect 82136 3760 135904 3788
rect 82136 3748 82142 3760
rect 135898 3748 135904 3760
rect 135956 3748 135962 3800
rect 209866 3748 209872 3800
rect 209924 3788 209930 3800
rect 229738 3788 229744 3800
rect 209924 3760 229744 3788
rect 209924 3748 209930 3760
rect 229738 3748 229744 3760
rect 229796 3748 229802 3800
rect 238110 3748 238116 3800
rect 238168 3788 238174 3800
rect 247678 3788 247684 3800
rect 238168 3760 247684 3788
rect 238168 3748 238174 3760
rect 247678 3748 247684 3760
rect 247736 3748 247742 3800
rect 318886 3748 318892 3800
rect 318944 3788 318950 3800
rect 330386 3788 330392 3800
rect 318944 3760 330392 3788
rect 318944 3748 318950 3760
rect 330386 3748 330392 3760
rect 330444 3748 330450 3800
rect 336734 3748 336740 3800
rect 336792 3788 336798 3800
rect 355226 3788 355232 3800
rect 336792 3760 355232 3788
rect 336792 3748 336798 3760
rect 355226 3748 355232 3760
rect 355284 3748 355290 3800
rect 390646 3748 390652 3800
rect 390704 3788 390710 3800
rect 433242 3788 433248 3800
rect 390704 3760 433248 3788
rect 390704 3748 390710 3760
rect 433242 3748 433248 3760
rect 433300 3748 433306 3800
rect 443638 3748 443644 3800
rect 443696 3788 443702 3800
rect 458082 3788 458088 3800
rect 443696 3760 458088 3788
rect 443696 3748 443702 3760
rect 458082 3748 458088 3760
rect 458140 3748 458146 3800
rect 478230 3748 478236 3800
rect 478288 3788 478294 3800
rect 539594 3788 539600 3800
rect 478288 3760 539600 3788
rect 478288 3748 478294 3760
rect 539594 3748 539600 3760
rect 539652 3748 539658 3800
rect 547138 3748 547144 3800
rect 547196 3788 547202 3800
rect 571518 3788 571524 3800
rect 547196 3760 571524 3788
rect 547196 3748 547202 3760
rect 571518 3748 571524 3760
rect 571576 3748 571582 3800
rect 46658 3680 46664 3732
rect 46716 3720 46722 3732
rect 117958 3720 117964 3732
rect 46716 3692 117964 3720
rect 46716 3680 46722 3692
rect 117958 3680 117964 3692
rect 118016 3680 118022 3732
rect 202690 3680 202696 3732
rect 202748 3720 202754 3732
rect 225598 3720 225604 3732
rect 202748 3692 225604 3720
rect 202748 3680 202754 3692
rect 225598 3680 225604 3692
rect 225656 3680 225662 3732
rect 234614 3680 234620 3732
rect 234672 3720 234678 3732
rect 246298 3720 246304 3732
rect 234672 3692 246304 3720
rect 234672 3680 234678 3692
rect 246298 3680 246304 3692
rect 246356 3680 246362 3732
rect 277118 3680 277124 3732
rect 277176 3720 277182 3732
rect 279418 3720 279424 3732
rect 277176 3692 279424 3720
rect 277176 3680 277182 3692
rect 279418 3680 279424 3692
rect 279476 3680 279482 3732
rect 279510 3680 279516 3732
rect 279568 3720 279574 3732
rect 283098 3720 283104 3732
rect 279568 3692 283104 3720
rect 279568 3680 279574 3692
rect 283098 3680 283104 3692
rect 283156 3680 283162 3732
rect 303706 3680 303712 3732
rect 303764 3720 303770 3732
rect 307938 3720 307944 3732
rect 303764 3692 307944 3720
rect 303764 3680 303770 3692
rect 307938 3680 307944 3692
rect 307996 3680 308002 3732
rect 320266 3680 320272 3732
rect 320324 3720 320330 3732
rect 332686 3720 332692 3732
rect 320324 3692 332692 3720
rect 320324 3680 320330 3692
rect 332686 3680 332692 3692
rect 332744 3680 332750 3732
rect 340874 3680 340880 3732
rect 340932 3720 340938 3732
rect 361114 3720 361120 3732
rect 340932 3692 361120 3720
rect 340932 3680 340938 3692
rect 361114 3680 361120 3692
rect 361172 3680 361178 3732
rect 362218 3680 362224 3732
rect 362276 3720 362282 3732
rect 372890 3720 372896 3732
rect 362276 3692 372896 3720
rect 362276 3680 362282 3692
rect 372890 3680 372896 3692
rect 372948 3680 372954 3732
rect 382918 3680 382924 3732
rect 382976 3720 382982 3732
rect 382976 3692 390692 3720
rect 382976 3680 382982 3692
rect 390664 3664 390692 3692
rect 391198 3680 391204 3732
rect 391256 3720 391262 3732
rect 394234 3720 394240 3732
rect 391256 3692 394240 3720
rect 391256 3680 391262 3692
rect 394234 3680 394240 3692
rect 394292 3680 394298 3732
rect 396074 3680 396080 3732
rect 396132 3720 396138 3732
rect 440326 3720 440332 3732
rect 396132 3692 440332 3720
rect 396132 3680 396138 3692
rect 440326 3680 440332 3692
rect 440384 3680 440390 3732
rect 446398 3680 446404 3732
rect 446456 3720 446462 3732
rect 461578 3720 461584 3732
rect 446456 3692 461584 3720
rect 446456 3680 446462 3692
rect 461578 3680 461584 3692
rect 461636 3680 461642 3732
rect 468478 3680 468484 3732
rect 468536 3720 468542 3732
rect 532510 3720 532516 3732
rect 468536 3692 532516 3720
rect 468536 3680 468542 3692
rect 532510 3680 532516 3692
rect 532568 3680 532574 3732
rect 548518 3680 548524 3732
rect 548576 3720 548582 3732
rect 578602 3720 578608 3732
rect 548576 3692 578608 3720
rect 548576 3680 548582 3692
rect 578602 3680 578608 3692
rect 578660 3680 578666 3732
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 114554 3652 114560 3664
rect 39632 3624 114560 3652
rect 39632 3612 39638 3624
rect 114554 3612 114560 3624
rect 114612 3612 114618 3664
rect 195606 3612 195612 3664
rect 195664 3652 195670 3664
rect 224218 3652 224224 3664
rect 195664 3624 224224 3652
rect 195664 3612 195670 3624
rect 224218 3612 224224 3624
rect 224276 3612 224282 3664
rect 231026 3612 231032 3664
rect 231084 3652 231090 3664
rect 242250 3652 242256 3664
rect 231084 3624 242256 3652
rect 231084 3612 231090 3624
rect 242250 3612 242256 3624
rect 242308 3612 242314 3664
rect 304994 3612 305000 3664
rect 305052 3652 305058 3664
rect 310238 3652 310244 3664
rect 305052 3624 310244 3652
rect 305052 3612 305058 3624
rect 310238 3612 310244 3624
rect 310296 3612 310302 3664
rect 313642 3612 313648 3664
rect 313700 3652 313706 3664
rect 323302 3652 323308 3664
rect 313700 3624 323308 3652
rect 313700 3612 313706 3624
rect 323302 3612 323308 3624
rect 323360 3612 323366 3664
rect 324590 3612 324596 3664
rect 324648 3652 324654 3664
rect 337470 3652 337476 3664
rect 324648 3624 337476 3652
rect 324648 3612 324654 3624
rect 337470 3612 337476 3624
rect 337528 3612 337534 3664
rect 338482 3612 338488 3664
rect 338540 3652 338546 3664
rect 358722 3652 358728 3664
rect 338540 3624 358728 3652
rect 338540 3612 338546 3624
rect 358722 3612 358728 3624
rect 358780 3612 358786 3664
rect 360838 3612 360844 3664
rect 360896 3652 360902 3664
rect 383562 3652 383568 3664
rect 360896 3624 383568 3652
rect 360896 3612 360902 3624
rect 383562 3612 383568 3624
rect 383620 3612 383626 3664
rect 390646 3612 390652 3664
rect 390704 3612 390710 3664
rect 400582 3612 400588 3664
rect 400640 3652 400646 3664
rect 447410 3652 447416 3664
rect 400640 3624 447416 3652
rect 400640 3612 400646 3624
rect 447410 3612 447416 3624
rect 447468 3612 447474 3664
rect 450538 3612 450544 3664
rect 450596 3652 450602 3664
rect 468662 3652 468668 3664
rect 450596 3624 468668 3652
rect 450596 3612 450602 3624
rect 468662 3612 468668 3624
rect 468720 3612 468726 3664
rect 472618 3612 472624 3664
rect 472676 3652 472682 3664
rect 546678 3652 546684 3664
rect 472676 3624 546684 3652
rect 472676 3612 472682 3624
rect 546678 3612 546684 3624
rect 546736 3612 546742 3664
rect 549898 3612 549904 3664
rect 549956 3652 549962 3664
rect 582190 3652 582196 3664
rect 549956 3624 582196 3652
rect 549956 3612 549962 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 10318 3584 10324 3596
rect 6886 3556 10324 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6886 3516 6914 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 98086 3584 98092 3596
rect 15988 3556 98092 3584
rect 15988 3544 15994 3556
rect 98086 3544 98092 3556
rect 98144 3544 98150 3596
rect 117590 3544 117596 3596
rect 117648 3584 117654 3596
rect 164878 3584 164884 3596
rect 117648 3556 164884 3584
rect 117648 3544 117654 3556
rect 164878 3544 164884 3556
rect 164936 3544 164942 3596
rect 181438 3544 181444 3596
rect 181496 3584 181502 3596
rect 181496 3556 188476 3584
rect 181496 3544 181502 3556
rect 5316 3488 6914 3516
rect 5316 3476 5322 3488
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 13078 3516 13084 3528
rect 10008 3488 13084 3516
rect 10008 3476 10014 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 97994 3516 98000 3528
rect 14792 3488 98000 3516
rect 14792 3476 14798 3488
rect 97994 3476 98000 3488
rect 98052 3476 98058 3528
rect 118694 3476 118700 3528
rect 118752 3516 118758 3528
rect 119890 3516 119896 3528
rect 118752 3488 119896 3516
rect 118752 3476 118758 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 121086 3476 121092 3528
rect 121144 3516 121150 3528
rect 167638 3516 167644 3528
rect 121144 3488 167644 3516
rect 121144 3476 121150 3488
rect 167638 3476 167644 3488
rect 167696 3476 167702 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 174630 3516 174636 3528
rect 173216 3488 174636 3516
rect 173216 3476 173222 3488
rect 174630 3476 174636 3488
rect 174688 3476 174694 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 178678 3516 178684 3528
rect 176712 3488 178684 3516
rect 176712 3476 176718 3488
rect 178678 3476 178684 3488
rect 178736 3476 178742 3528
rect 187326 3476 187332 3528
rect 187384 3516 187390 3528
rect 188338 3516 188344 3528
rect 187384 3488 188344 3516
rect 187384 3476 187390 3488
rect 188338 3476 188344 3488
rect 188396 3476 188402 3528
rect 188448 3516 188476 3556
rect 188522 3544 188528 3596
rect 188580 3584 188586 3596
rect 219526 3584 219532 3596
rect 188580 3556 219532 3584
rect 188580 3544 188586 3556
rect 219526 3544 219532 3556
rect 219584 3544 219590 3596
rect 227530 3544 227536 3596
rect 227588 3584 227594 3596
rect 239398 3584 239404 3596
rect 227588 3556 239404 3584
rect 227588 3544 227594 3556
rect 239398 3544 239404 3556
rect 239456 3544 239462 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 252370 3584 252376 3596
rect 251232 3556 252376 3584
rect 251232 3544 251238 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 258258 3544 258264 3596
rect 258316 3584 258322 3596
rect 261478 3584 261484 3596
rect 258316 3556 261484 3584
rect 258316 3544 258322 3556
rect 261478 3544 261484 3556
rect 261536 3544 261542 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 268470 3584 268476 3596
rect 267792 3556 268476 3584
rect 267792 3544 267798 3556
rect 268470 3544 268476 3556
rect 268528 3544 268534 3596
rect 283098 3544 283104 3596
rect 283156 3584 283162 3596
rect 285766 3584 285772 3596
rect 283156 3556 285772 3584
rect 283156 3544 283162 3556
rect 285766 3544 285772 3556
rect 285824 3544 285830 3596
rect 317782 3544 317788 3596
rect 317840 3584 317846 3596
rect 329190 3584 329196 3596
rect 317840 3556 329196 3584
rect 317840 3544 317846 3556
rect 329190 3544 329196 3556
rect 329248 3544 329254 3596
rect 331306 3544 331312 3596
rect 331364 3584 331370 3596
rect 348050 3584 348056 3596
rect 331364 3556 348056 3584
rect 331364 3544 331370 3556
rect 348050 3544 348056 3556
rect 348108 3544 348114 3596
rect 350902 3544 350908 3596
rect 350960 3584 350966 3596
rect 376478 3584 376484 3596
rect 350960 3556 376484 3584
rect 350960 3544 350966 3556
rect 376478 3544 376484 3556
rect 376536 3544 376542 3596
rect 377398 3544 377404 3596
rect 377456 3584 377462 3596
rect 387150 3584 387156 3596
rect 377456 3556 387156 3584
rect 377456 3544 377462 3556
rect 387150 3544 387156 3556
rect 387208 3544 387214 3596
rect 405734 3544 405740 3596
rect 405792 3584 405798 3596
rect 454494 3584 454500 3596
rect 405792 3556 454500 3584
rect 405792 3544 405798 3556
rect 454494 3544 454500 3556
rect 454552 3544 454558 3596
rect 482278 3544 482284 3596
rect 482336 3584 482342 3596
rect 560846 3584 560852 3596
rect 482336 3556 560852 3584
rect 482336 3544 482342 3556
rect 560846 3544 560852 3556
rect 560904 3544 560910 3596
rect 213914 3516 213920 3528
rect 188448 3488 213920 3516
rect 213914 3476 213920 3488
rect 213972 3476 213978 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 228358 3516 228364 3528
rect 226392 3488 228364 3516
rect 226392 3476 226398 3488
rect 228358 3476 228364 3488
rect 228416 3476 228422 3528
rect 242158 3516 242164 3528
rect 228560 3488 242164 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 92474 3448 92480 3460
rect 6512 3420 92480 3448
rect 6512 3408 6518 3420
rect 92474 3408 92480 3420
rect 92532 3408 92538 3460
rect 96246 3408 96252 3460
rect 96304 3448 96310 3460
rect 144178 3448 144184 3460
rect 96304 3420 144184 3448
rect 96304 3408 96310 3420
rect 144178 3408 144184 3420
rect 144236 3408 144242 3460
rect 160094 3408 160100 3460
rect 160152 3448 160158 3460
rect 160152 3420 161474 3448
rect 160152 3408 160158 3420
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 32398 3380 32404 3392
rect 28960 3352 32404 3380
rect 28960 3340 28966 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 69014 3340 69020 3392
rect 69072 3380 69078 3392
rect 69934 3380 69940 3392
rect 69072 3352 69940 3380
rect 69072 3340 69078 3352
rect 69934 3340 69940 3352
rect 69992 3340 69998 3392
rect 161446 3380 161474 3420
rect 174262 3408 174268 3460
rect 174320 3448 174326 3460
rect 175918 3448 175924 3460
rect 174320 3420 175924 3448
rect 174320 3408 174326 3420
rect 175918 3408 175924 3420
rect 175976 3408 175982 3460
rect 177850 3408 177856 3460
rect 177908 3448 177914 3460
rect 210418 3448 210424 3460
rect 177908 3420 210424 3448
rect 177908 3408 177914 3420
rect 210418 3408 210424 3420
rect 210476 3408 210482 3460
rect 219250 3408 219256 3460
rect 219308 3448 219314 3460
rect 219308 3420 219434 3448
rect 219308 3408 219314 3420
rect 174538 3380 174544 3392
rect 161446 3352 174544 3380
rect 174538 3340 174544 3352
rect 174596 3340 174602 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 192478 3380 192484 3392
rect 190880 3352 192484 3380
rect 190880 3340 190886 3352
rect 192478 3340 192484 3352
rect 192536 3340 192542 3392
rect 209774 3340 209780 3392
rect 209832 3380 209838 3392
rect 210970 3380 210976 3392
rect 209832 3352 210976 3380
rect 209832 3340 209838 3352
rect 210970 3340 210976 3352
rect 211028 3340 211034 3392
rect 2866 3272 2872 3324
rect 2924 3312 2930 3324
rect 8938 3312 8944 3324
rect 2924 3284 8944 3312
rect 2924 3272 2930 3284
rect 8938 3272 8944 3284
rect 8996 3272 9002 3324
rect 19426 3272 19432 3324
rect 19484 3312 19490 3324
rect 25498 3312 25504 3324
rect 19484 3284 25504 3312
rect 19484 3272 19490 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 219406 3312 219434 3420
rect 222746 3340 222752 3392
rect 222804 3380 222810 3392
rect 228560 3380 228588 3488
rect 242158 3476 242164 3488
rect 242216 3476 242222 3528
rect 245194 3476 245200 3528
rect 245252 3516 245258 3528
rect 255958 3516 255964 3528
rect 245252 3488 255964 3516
rect 245252 3476 245258 3488
rect 255958 3476 255964 3488
rect 256016 3476 256022 3528
rect 272426 3476 272432 3528
rect 272484 3516 272490 3528
rect 273898 3516 273904 3528
rect 272484 3488 273904 3516
rect 272484 3476 272490 3488
rect 273898 3476 273904 3488
rect 273956 3476 273962 3528
rect 300946 3476 300952 3528
rect 301004 3516 301010 3528
rect 305546 3516 305552 3528
rect 301004 3488 305552 3516
rect 301004 3476 301010 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 313826 3516 313832 3528
rect 309836 3488 313832 3516
rect 309836 3476 309842 3488
rect 313826 3476 313832 3488
rect 313884 3476 313890 3528
rect 323026 3476 323032 3528
rect 323084 3516 323090 3528
rect 336274 3516 336280 3528
rect 323084 3488 336280 3516
rect 323084 3476 323090 3488
rect 336274 3476 336280 3488
rect 336332 3476 336338 3528
rect 341058 3476 341064 3528
rect 341116 3516 341122 3528
rect 362310 3516 362316 3528
rect 341116 3488 362316 3516
rect 341116 3476 341122 3488
rect 362310 3476 362316 3488
rect 362368 3476 362374 3528
rect 369118 3476 369124 3528
rect 369176 3516 369182 3528
rect 397730 3516 397736 3528
rect 369176 3488 397736 3516
rect 369176 3476 369182 3488
rect 397730 3476 397736 3488
rect 397788 3476 397794 3528
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 400858 3476 400864 3528
rect 400916 3516 400922 3528
rect 411898 3516 411904 3528
rect 400916 3488 411904 3516
rect 400916 3476 400922 3488
rect 411898 3476 411904 3488
rect 411956 3476 411962 3528
rect 412634 3476 412640 3528
rect 412692 3516 412698 3528
rect 465166 3516 465172 3528
rect 412692 3488 465172 3516
rect 412692 3476 412698 3488
rect 465166 3476 465172 3488
rect 465224 3476 465230 3528
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474182 3516 474188 3528
rect 473412 3488 474188 3516
rect 473412 3476 473418 3488
rect 474182 3476 474188 3488
rect 474240 3476 474246 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 494054 3476 494060 3528
rect 494112 3516 494118 3528
rect 580994 3516 581000 3528
rect 494112 3488 581000 3516
rect 494112 3476 494118 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 238018 3448 238024 3460
rect 222804 3352 228588 3380
rect 229066 3420 238024 3448
rect 222804 3340 222810 3352
rect 229066 3312 229094 3420
rect 238018 3408 238024 3420
rect 238076 3408 238082 3460
rect 240502 3408 240508 3460
rect 240560 3448 240566 3460
rect 253198 3448 253204 3460
rect 240560 3420 253204 3448
rect 240560 3408 240566 3420
rect 253198 3408 253204 3420
rect 253256 3408 253262 3460
rect 290182 3408 290188 3460
rect 290240 3448 290246 3460
rect 291194 3448 291200 3460
rect 290240 3420 291200 3448
rect 290240 3408 290246 3420
rect 291194 3408 291200 3420
rect 291252 3408 291258 3460
rect 296806 3408 296812 3460
rect 296864 3448 296870 3460
rect 299658 3448 299664 3460
rect 296864 3420 299664 3448
rect 296864 3408 296870 3420
rect 299658 3408 299664 3420
rect 299716 3408 299722 3460
rect 307018 3408 307024 3460
rect 307076 3448 307082 3460
rect 311434 3448 311440 3460
rect 307076 3420 311440 3448
rect 307076 3408 307082 3420
rect 311434 3408 311440 3420
rect 311492 3408 311498 3460
rect 313366 3408 313372 3460
rect 313424 3448 313430 3460
rect 322106 3448 322112 3460
rect 313424 3420 322112 3448
rect 313424 3408 313430 3420
rect 322106 3408 322112 3420
rect 322164 3408 322170 3460
rect 326062 3408 326068 3460
rect 326120 3448 326126 3460
rect 340966 3448 340972 3460
rect 326120 3420 340972 3448
rect 326120 3408 326126 3420
rect 340966 3408 340972 3420
rect 341024 3408 341030 3460
rect 349154 3408 349160 3460
rect 349212 3448 349218 3460
rect 350442 3448 350448 3460
rect 349212 3420 350448 3448
rect 349212 3408 349218 3420
rect 350442 3408 350448 3420
rect 350500 3408 350506 3460
rect 369394 3448 369400 3460
rect 354646 3420 369400 3448
rect 310514 3340 310520 3392
rect 310572 3380 310578 3392
rect 318518 3380 318524 3392
rect 310572 3352 318524 3380
rect 310572 3340 310578 3352
rect 318518 3340 318524 3352
rect 318576 3340 318582 3392
rect 346578 3340 346584 3392
rect 346636 3380 346642 3392
rect 354646 3380 354674 3420
rect 369394 3408 369400 3420
rect 369452 3408 369458 3460
rect 371234 3408 371240 3460
rect 371292 3448 371298 3460
rect 404814 3448 404820 3460
rect 371292 3420 404820 3448
rect 371292 3408 371298 3420
rect 404814 3408 404820 3420
rect 404872 3408 404878 3460
rect 418246 3408 418252 3460
rect 418304 3448 418310 3460
rect 472250 3448 472256 3460
rect 418304 3420 472256 3448
rect 418304 3408 418310 3420
rect 472250 3408 472256 3420
rect 472308 3408 472314 3460
rect 495526 3408 495532 3460
rect 495584 3448 495590 3460
rect 583386 3448 583392 3460
rect 495584 3420 583392 3448
rect 495584 3408 495590 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 346636 3352 354674 3380
rect 346636 3340 346642 3352
rect 435358 3340 435364 3392
rect 435416 3380 435422 3392
rect 436738 3380 436744 3392
rect 435416 3352 436744 3380
rect 435416 3340 435422 3352
rect 436738 3340 436744 3352
rect 436796 3340 436802 3392
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 548702 3380 548708 3392
rect 547932 3352 548708 3380
rect 547932 3340 547938 3352
rect 548702 3340 548708 3352
rect 548760 3340 548766 3392
rect 219406 3284 229094 3312
rect 311158 3272 311164 3324
rect 311216 3312 311222 3324
rect 315022 3312 315028 3324
rect 311216 3284 315028 3312
rect 311216 3272 311222 3284
rect 315022 3272 315028 3284
rect 315080 3272 315086 3324
rect 318058 3272 318064 3324
rect 318116 3312 318122 3324
rect 325602 3312 325608 3324
rect 318116 3284 325608 3312
rect 318116 3272 318122 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 358078 3272 358084 3324
rect 358136 3312 358142 3324
rect 365806 3312 365812 3324
rect 358136 3284 365812 3312
rect 358136 3272 358142 3284
rect 365806 3272 365812 3284
rect 365864 3272 365870 3324
rect 374638 3272 374644 3324
rect 374696 3312 374702 3324
rect 379974 3312 379980 3324
rect 374696 3284 379980 3312
rect 374696 3272 374702 3284
rect 379974 3272 379980 3284
rect 380032 3272 380038 3324
rect 11146 3204 11152 3256
rect 11204 3244 11210 3256
rect 14458 3244 14464 3256
rect 11204 3216 14464 3244
rect 11204 3204 11210 3216
rect 14458 3204 14464 3216
rect 14516 3204 14522 3256
rect 309318 3204 309324 3256
rect 309376 3244 309382 3256
rect 316218 3244 316224 3256
rect 309376 3216 316224 3244
rect 309376 3204 309382 3216
rect 316218 3204 316224 3216
rect 316276 3204 316282 3256
rect 576118 3204 576124 3256
rect 576176 3244 576182 3256
rect 577406 3244 577412 3256
rect 576176 3216 577412 3244
rect 576176 3204 576182 3216
rect 577406 3204 577412 3216
rect 577464 3204 577470 3256
rect 35986 3136 35992 3188
rect 36044 3176 36050 3188
rect 39298 3176 39304 3188
rect 36044 3148 39304 3176
rect 36044 3136 36050 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 167178 3136 167184 3188
rect 167236 3176 167242 3188
rect 170398 3176 170404 3188
rect 167236 3148 170404 3176
rect 167236 3136 167242 3148
rect 170398 3136 170404 3148
rect 170456 3136 170462 3188
rect 540238 3136 540244 3188
rect 540296 3176 540302 3188
rect 543182 3176 543188 3188
rect 540296 3148 543188 3176
rect 540296 3136 540302 3148
rect 543182 3136 543188 3148
rect 543240 3136 543246 3188
rect 566 3068 572 3120
rect 624 3108 630 3120
rect 4798 3108 4804 3120
rect 624 3080 4804 3108
rect 624 3068 630 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 309134 3068 309140 3120
rect 309192 3108 309198 3120
rect 317322 3108 317328 3120
rect 309192 3080 317328 3108
rect 309192 3068 309198 3080
rect 317322 3068 317328 3080
rect 317380 3068 317386 3120
rect 155402 3000 155408 3052
rect 155460 3040 155466 3052
rect 157978 3040 157984 3052
rect 155460 3012 157984 3040
rect 155460 3000 155466 3012
rect 157978 3000 157984 3012
rect 158036 3000 158042 3052
rect 295426 3000 295432 3052
rect 295484 3040 295490 3052
rect 297266 3040 297272 3052
rect 295484 3012 297272 3040
rect 295484 3000 295490 3012
rect 297266 3000 297272 3012
rect 297324 3000 297330 3052
rect 303522 3000 303528 3052
rect 303580 3040 303586 3052
rect 306742 3040 306748 3052
rect 303580 3012 306748 3040
rect 303580 3000 303586 3012
rect 306742 3000 306748 3012
rect 306800 3000 306806 3052
rect 296898 2932 296904 2984
rect 296956 2972 296962 2984
rect 298462 2972 298468 2984
rect 296956 2944 298468 2972
rect 296956 2932 296962 2944
rect 298462 2932 298468 2944
rect 298520 2932 298526 2984
rect 306466 2932 306472 2984
rect 306524 2972 306530 2984
rect 312630 2972 312636 2984
rect 306524 2944 312636 2972
rect 306524 2932 306530 2944
rect 312630 2932 312636 2944
rect 312688 2932 312694 2984
rect 393958 2932 393964 2984
rect 394016 2972 394022 2984
rect 401318 2972 401324 2984
rect 394016 2944 401324 2972
rect 394016 2932 394022 2944
rect 401318 2932 401324 2944
rect 401376 2932 401382 2984
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 283840 700884 283892 700936
rect 301412 700884 301464 700936
rect 290096 700816 290148 700868
rect 348792 700816 348844 700868
rect 218980 700748 219032 700800
rect 312728 700748 312780 700800
rect 278780 700680 278832 700732
rect 413652 700680 413704 700732
rect 154120 700612 154172 700664
rect 324044 700612 324096 700664
rect 267464 700544 267516 700596
rect 478512 700544 478564 700596
rect 89168 700476 89220 700528
rect 335360 700476 335412 700528
rect 256148 700408 256200 700460
rect 543464 700408 543516 700460
rect 24308 700340 24360 700392
rect 346676 700340 346728 700392
rect 8116 700272 8168 700324
rect 342904 700272 342956 700324
rect 549904 700272 549956 700324
rect 559656 700272 559708 700324
rect 267648 698980 267700 699032
rect 297640 698980 297692 699032
rect 275008 698912 275060 698964
rect 397460 698912 397512 698964
rect 137836 697552 137888 697604
rect 320272 697552 320324 697604
rect 241060 696940 241112 696992
rect 580172 696940 580224 696992
rect 105452 696192 105504 696244
rect 327816 696192 327868 696244
rect 244832 683204 244884 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 350448 683136 350500 683188
rect 237288 670760 237340 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 357992 670692 358044 670744
rect 286324 663008 286376 663060
rect 331220 663008 331272 663060
rect 3424 656888 3476 656940
rect 354220 656888 354272 656940
rect 229744 643084 229796 643136
rect 580172 643084 580224 643136
rect 201500 642336 201552 642388
rect 308956 642336 309008 642388
rect 234620 640976 234672 641028
rect 305184 640976 305236 641028
rect 263692 639548 263744 639600
rect 462320 639548 462372 639600
rect 71780 638392 71832 638444
rect 331588 638392 331640 638444
rect 252376 638324 252428 638376
rect 527180 638324 527232 638376
rect 68376 638256 68428 638308
rect 369308 638256 369360 638308
rect 184480 638188 184532 638240
rect 522396 638188 522448 638240
rect 58624 638120 58676 638172
rect 403256 638120 403308 638172
rect 173164 638052 173216 638104
rect 521016 638052 521068 638104
rect 161848 637984 161900 638036
rect 520924 637984 520976 638036
rect 57244 637916 57296 637968
rect 422116 637916 422168 637968
rect 150532 637848 150584 637900
rect 518256 637848 518308 637900
rect 7564 637780 7616 637832
rect 388168 637780 388220 637832
rect 13084 637712 13136 637764
rect 410432 637712 410484 637764
rect 109040 637644 109092 637696
rect 515404 637644 515456 637696
rect 105268 637576 105320 637628
rect 516784 637576 516836 637628
rect 169760 637100 169812 637152
rect 316132 637100 316184 637152
rect 40040 637032 40092 637084
rect 338764 637032 338816 637084
rect 248880 636964 248932 637016
rect 549904 636964 549956 637016
rect 180708 636896 180760 636948
rect 516968 636896 517020 636948
rect 53104 636828 53156 636880
rect 414204 636828 414256 636880
rect 147036 636760 147088 636812
rect 516876 636760 516928 636812
rect 66904 636692 66956 636744
rect 440608 636692 440660 636744
rect 124128 636624 124180 636676
rect 514208 636624 514260 636676
rect 71044 636556 71096 636608
rect 463240 636556 463292 636608
rect 64144 636488 64196 636540
rect 474740 636488 474792 636540
rect 68284 636420 68336 636472
rect 485872 636420 485924 636472
rect 72424 636352 72476 636404
rect 497188 636352 497240 636404
rect 21364 636284 21416 636336
rect 451924 636284 451976 636336
rect 94228 636216 94280 636268
rect 531964 636216 532016 636268
rect 293868 635672 293920 635724
rect 299480 635672 299532 635724
rect 282828 635604 282880 635656
rect 364340 635604 364392 635656
rect 271512 635536 271564 635588
rect 429200 635536 429252 635588
rect 260196 635468 260248 635520
rect 494060 635468 494112 635520
rect 226248 635400 226300 635452
rect 512828 635400 512880 635452
rect 214932 635332 214984 635384
rect 512736 635332 512788 635384
rect 71320 635264 71372 635316
rect 372712 635264 372764 635316
rect 203616 635196 203668 635248
rect 514300 635196 514352 635248
rect 71228 635128 71280 635180
rect 384028 635128 384080 635180
rect 199844 635060 199896 635112
rect 525248 635060 525300 635112
rect 62764 634992 62816 635044
rect 395344 634992 395396 635044
rect 71136 634924 71188 634976
rect 406660 634924 406712 634976
rect 3516 634856 3568 634908
rect 361580 634856 361632 634908
rect 113088 634788 113140 634840
rect 514116 634788 514168 634840
rect 216680 634312 216732 634364
rect 433432 634312 433484 634364
rect 139308 634244 139360 634296
rect 365628 634244 365680 634296
rect 366548 634244 366600 634296
rect 459560 634244 459612 634296
rect 177212 634176 177264 634228
rect 525156 634176 525208 634228
rect 192300 634108 192352 634160
rect 545764 634108 545816 634160
rect 165896 634040 165948 634092
rect 525064 634040 525116 634092
rect 154488 633972 154540 634024
rect 522304 633972 522356 634024
rect 131948 633904 132000 633956
rect 518164 633904 518216 633956
rect 4068 633836 4120 633888
rect 391940 633836 391992 633888
rect 3884 633768 3936 633820
rect 425520 633768 425572 633820
rect 3792 633700 3844 633752
rect 436836 633700 436888 633752
rect 4988 633632 5040 633684
rect 448520 633632 448572 633684
rect 3424 633564 3476 633616
rect 455696 633564 455748 633616
rect 505376 633564 505428 633616
rect 512000 633564 512052 633616
rect 4896 633496 4948 633548
rect 470876 633496 470928 633548
rect 501604 633496 501656 633548
rect 511080 633496 511132 633548
rect 4804 633428 4856 633480
rect 482100 633428 482152 633480
rect 493968 633428 494020 633480
rect 512092 633428 512144 633480
rect 5264 632884 5316 632936
rect 365168 632884 365220 632936
rect 158352 632816 158404 632868
rect 511448 632816 511500 632868
rect 3700 632748 3752 632800
rect 216680 632748 216732 632800
rect 222476 632748 222528 632800
rect 579988 632748 580040 632800
rect 365628 632680 365680 632732
rect 580448 632680 580500 632732
rect 218704 632612 218756 632664
rect 580080 632612 580132 632664
rect 3332 632544 3384 632596
rect 376852 632544 376904 632596
rect 207388 632476 207440 632528
rect 580908 632476 580960 632528
rect 135720 632408 135772 632460
rect 511356 632408 511408 632460
rect 3240 632340 3292 632392
rect 380256 632340 380308 632392
rect 195888 632272 195940 632324
rect 580724 632272 580776 632324
rect 3976 632204 4028 632256
rect 399116 632204 399168 632256
rect 3608 632136 3660 632188
rect 444702 632136 444754 632188
rect 127854 632068 127906 632120
rect 580264 632068 580316 632120
rect 410064 631660 410116 631712
rect 421012 631660 421064 631712
rect 142804 631524 142856 631576
rect 146944 631524 146996 631576
rect 5172 630776 5224 630828
rect 5080 630708 5132 630760
rect 142804 631388 142856 631440
rect 143264 631388 143316 631440
rect 146944 631388 146996 631440
rect 169668 631388 169720 631440
rect 188528 631388 188580 631440
rect 211068 631388 211120 631440
rect 233792 631388 233844 631440
rect 410064 631388 410116 631440
rect 410524 631388 410576 631440
rect 415492 631388 415544 631440
rect 421012 631456 421064 631508
rect 416596 631388 416648 631440
rect 429292 631388 429344 631440
rect 580172 631048 580224 631100
rect 580816 630980 580868 631032
rect 580632 630912 580684 630964
rect 580540 630844 580592 630896
rect 579988 630708 580040 630760
rect 580172 630708 580224 630760
rect 580356 630640 580408 630692
rect 3148 619556 3200 619608
rect 68376 619556 68428 619608
rect 512828 618196 512880 618248
rect 579988 618196 580040 618248
rect 2780 607044 2832 607096
rect 5264 607044 5316 607096
rect 3148 580932 3200 580984
rect 71320 580932 71372 580984
rect 512736 564340 512788 564392
rect 580172 564340 580224 564392
rect 3332 528504 3384 528556
rect 71228 528504 71280 528556
rect 514300 511912 514352 511964
rect 580172 511912 580224 511964
rect 3332 501780 3384 501832
rect 7564 501780 7616 501832
rect 3332 476008 3384 476060
rect 62764 476008 62816 476060
rect 525248 471928 525300 471980
rect 579804 471928 579856 471980
rect 3332 463632 3384 463684
rect 58624 463632 58676 463684
rect 545764 458124 545816 458176
rect 580172 458124 580224 458176
rect 522396 431876 522448 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 71136 423580 71188 423632
rect 3332 411204 3384 411256
rect 53104 411204 53156 411256
rect 516968 405628 517020 405680
rect 580172 405628 580224 405680
rect 3332 398760 3384 398812
rect 13084 398760 13136 398812
rect 521016 379448 521068 379500
rect 579620 379448 579672 379500
rect 2780 372308 2832 372360
rect 5172 372308 5224 372360
rect 525156 365644 525208 365696
rect 580172 365644 580224 365696
rect 2964 346332 3016 346384
rect 57244 346332 57296 346384
rect 520924 325592 520976 325644
rect 580172 325592 580224 325644
rect 2780 319812 2832 319864
rect 5080 319812 5132 319864
rect 525064 313216 525116 313268
rect 579712 313216 579764 313268
rect 511448 299412 511500 299464
rect 579804 299412 579856 299464
rect 518256 273164 518308 273216
rect 580172 273164 580224 273216
rect 3240 267656 3292 267708
rect 66904 267656 66956 267708
rect 522304 259360 522356 259412
rect 580172 259360 580224 259412
rect 2780 254940 2832 254992
rect 4988 254940 5040 254992
rect 516876 245556 516928 245608
rect 580172 245556 580224 245608
rect 3332 215228 3384 215280
rect 21364 215228 21416 215280
rect 511356 206932 511408 206984
rect 580172 206932 580224 206984
rect 518164 179324 518216 179376
rect 580172 179324 580224 179376
rect 514208 166948 514260 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 71044 164160 71096 164212
rect 2780 149880 2832 149932
rect 4896 149880 4948 149932
rect 514116 126896 514168 126948
rect 580172 126896 580224 126948
rect 516784 113092 516836 113144
rect 579804 113092 579856 113144
rect 3424 111732 3476 111784
rect 64144 111732 64196 111784
rect 515404 100648 515456 100700
rect 580172 100648 580224 100700
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 511264 86912 511316 86964
rect 580172 86912 580224 86964
rect 531964 73108 532016 73160
rect 580172 73108 580224 73160
rect 89720 71884 89772 71936
rect 90778 71884 90830 71936
rect 110420 71884 110472 71936
rect 111478 71884 111530 71936
rect 114560 71884 114612 71936
rect 115618 71884 115670 71936
rect 122840 71884 122892 71936
rect 123898 71884 123950 71936
rect 131120 71884 131172 71936
rect 132178 71884 132230 71936
rect 135260 71884 135312 71936
rect 136318 71884 136370 71936
rect 147680 71884 147732 71936
rect 148738 71884 148790 71936
rect 160100 71884 160152 71936
rect 161158 71884 161210 71936
rect 176660 71884 176712 71936
rect 177718 71884 177770 71936
rect 197452 71884 197504 71936
rect 198418 71884 198470 71936
rect 201500 71884 201552 71936
rect 202558 71884 202610 71936
rect 213920 71884 213972 71936
rect 214978 71884 215030 71936
rect 296812 71884 296864 71936
rect 297778 71884 297830 71936
rect 309140 71884 309192 71936
rect 310198 71884 310250 71936
rect 346492 71884 346544 71936
rect 347458 71884 347510 71936
rect 367100 71884 367152 71936
rect 368158 71884 368210 71936
rect 412640 71884 412692 71936
rect 413698 71884 413750 71936
rect 441620 71884 441672 71936
rect 442678 71884 442730 71936
rect 3424 71680 3476 71732
rect 68284 71680 68336 71732
rect 233332 70320 233384 70372
rect 251364 70320 251416 70372
rect 246304 70252 246356 70304
rect 252192 70252 252244 70304
rect 77300 70184 77352 70236
rect 142896 70184 142948 70236
rect 238024 70184 238076 70236
rect 241520 70184 241572 70236
rect 247684 70184 247736 70236
rect 254676 70184 254728 70236
rect 260840 70184 260892 70236
rect 271236 70184 271288 70236
rect 50344 70116 50396 70168
rect 118056 70116 118108 70168
rect 217324 70116 217376 70168
rect 229100 70116 229152 70168
rect 256700 70116 256752 70168
rect 267924 70116 267976 70168
rect 483296 70116 483348 70168
rect 494704 70184 494756 70236
rect 494888 70184 494940 70236
rect 549904 70184 549956 70236
rect 493232 70116 493284 70168
rect 548524 70116 548576 70168
rect 70400 70048 70452 70100
rect 138020 70048 138072 70100
rect 198740 70048 198792 70100
rect 227352 70048 227404 70100
rect 254032 70048 254084 70100
rect 266360 70048 266412 70100
rect 359096 70048 359148 70100
rect 377404 70048 377456 70100
rect 416228 70048 416280 70100
rect 450544 70048 450596 70100
rect 488264 70048 488316 70100
rect 39304 69980 39356 70032
rect 113180 69980 113232 70032
rect 174544 69980 174596 70032
rect 200120 69980 200172 70032
rect 221464 69980 221516 70032
rect 233976 69980 234028 70032
rect 248420 69980 248472 70032
rect 262220 69980 262272 70032
rect 263600 69980 263652 70032
rect 272892 69980 272944 70032
rect 273260 69980 273312 70032
rect 279516 69980 279568 70032
rect 361580 69980 361632 70032
rect 382924 69980 382976 70032
rect 408776 69980 408828 70032
rect 443644 69980 443696 70032
rect 465908 69980 465960 70032
rect 478144 69980 478196 70032
rect 547144 70048 547196 70100
rect 494704 69980 494756 70032
rect 545764 69980 545816 70032
rect 28264 69912 28316 69964
rect 102324 69912 102376 69964
rect 135904 69912 135956 69964
rect 145380 69912 145432 69964
rect 197360 69912 197412 69964
rect 226524 69912 226576 69964
rect 228364 69912 228416 69964
rect 246396 69912 246448 69964
rect 247040 69912 247092 69964
rect 261300 69912 261352 69964
rect 266360 69912 266412 69964
rect 274640 69912 274692 69964
rect 320180 69912 320232 69964
rect 327724 69912 327776 69964
rect 374000 69912 374052 69964
rect 398104 69912 398156 69964
rect 421196 69912 421248 69964
rect 474740 69912 474792 69964
rect 478328 69912 478380 69964
rect 543004 69912 543056 69964
rect 32404 69844 32456 69896
rect 108120 69844 108172 69896
rect 140044 69844 140096 69896
rect 150440 69844 150492 69896
rect 167644 69844 167696 69896
rect 172520 69844 172572 69896
rect 191840 69844 191892 69896
rect 222384 69844 222436 69896
rect 225604 69844 225656 69896
rect 229836 69844 229888 69896
rect 235264 69844 235316 69896
rect 239772 69844 239824 69896
rect 251272 69844 251324 69896
rect 263784 69844 263836 69896
rect 264980 69844 265032 69896
rect 273720 69844 273772 69896
rect 273904 69844 273956 69896
rect 278780 69844 278832 69896
rect 306104 69844 306156 69896
rect 307024 69844 307076 69896
rect 334256 69844 334308 69896
rect 336004 69844 336056 69896
rect 350816 69844 350868 69896
rect 355324 69844 355376 69896
rect 25504 69776 25556 69828
rect 101496 69776 101548 69828
rect 144184 69776 144236 69828
rect 155316 69776 155368 69828
rect 156604 69776 156656 69828
rect 167736 69776 167788 69828
rect 170404 69776 170456 69828
rect 204996 69776 205048 69828
rect 205640 69776 205692 69828
rect 232320 69776 232372 69828
rect 236000 69776 236052 69828
rect 253940 69776 253992 69828
rect 255320 69776 255372 69828
rect 267096 69776 267148 69828
rect 285680 69776 285732 69828
rect 288624 69776 288676 69828
rect 354128 69776 354180 69828
rect 374644 69844 374696 69896
rect 376484 69844 376536 69896
rect 400864 69844 400916 69896
rect 411260 69844 411312 69896
rect 446404 69844 446456 69896
rect 453488 69844 453540 69896
rect 521660 69844 521712 69896
rect 369032 69776 369084 69828
rect 393964 69776 394016 69828
rect 403808 69776 403860 69828
rect 440884 69776 440936 69828
rect 445760 69776 445812 69828
rect 453304 69776 453356 69828
rect 458456 69776 458508 69828
rect 528560 69776 528612 69828
rect 14464 69708 14516 69760
rect 95700 69708 95752 69760
rect 124220 69708 124272 69760
rect 175280 69708 175332 69760
rect 184940 69708 184992 69760
rect 217416 69708 217468 69760
rect 229100 69708 229152 69760
rect 248880 69708 248932 69760
rect 251180 69708 251232 69760
rect 264612 69708 264664 69760
rect 335912 69708 335964 69760
rect 345664 69708 345716 69760
rect 349160 69708 349212 69760
rect 362224 69708 362276 69760
rect 10324 69640 10376 69692
rect 91560 69640 91612 69692
rect 106280 69640 106332 69692
rect 162860 69640 162912 69692
rect 169760 69640 169812 69692
rect 207480 69640 207532 69692
rect 219440 69640 219492 69692
rect 242256 69640 242308 69692
rect 242900 69640 242952 69692
rect 258816 69640 258868 69692
rect 259460 69640 259512 69692
rect 270500 69640 270552 69692
rect 274640 69640 274692 69692
rect 280344 69640 280396 69692
rect 311900 69640 311952 69692
rect 318800 69640 318852 69692
rect 325976 69640 326028 69692
rect 336096 69640 336148 69692
rect 344192 69640 344244 69692
rect 358084 69640 358136 69692
rect 358268 69640 358320 69692
rect 385040 69708 385092 69760
rect 398840 69708 398892 69760
rect 436744 69708 436796 69760
rect 468392 69708 468444 69760
rect 540244 69708 540296 69760
rect 364064 69640 364116 69692
rect 391204 69640 391256 69692
rect 393872 69640 393924 69692
rect 435364 69640 435416 69692
rect 448520 69640 448572 69692
rect 456064 69640 456116 69692
rect 463424 69640 463476 69692
rect 535460 69640 535512 69692
rect 233884 69504 233936 69556
rect 238944 69504 238996 69556
rect 242256 69504 242308 69556
rect 249800 69504 249852 69556
rect 270500 69504 270552 69556
rect 277860 69504 277912 69556
rect 267740 69300 267792 69352
rect 276204 69300 276256 69352
rect 261484 69232 261536 69284
rect 268752 69232 268804 69284
rect 277400 69232 277452 69284
rect 282920 69232 282972 69284
rect 284300 69232 284352 69284
rect 287796 69232 287848 69284
rect 300860 69232 300912 69284
rect 303620 69232 303672 69284
rect 267832 69164 267884 69216
rect 275376 69164 275428 69216
rect 280160 69164 280212 69216
rect 284484 69164 284536 69216
rect 164884 69096 164936 69148
rect 170220 69096 170272 69148
rect 239404 69096 239456 69148
rect 247224 69096 247276 69148
rect 269120 69096 269172 69148
rect 277032 69096 277084 69148
rect 278044 69096 278096 69148
rect 281172 69096 281224 69148
rect 281540 69096 281592 69148
rect 285312 69096 285364 69148
rect 287060 69096 287112 69148
rect 289452 69096 289504 69148
rect 299480 69096 299532 69148
rect 300860 69096 300912 69148
rect 308588 69096 308640 69148
rect 311164 69096 311216 69148
rect 317696 69096 317748 69148
rect 323584 69096 323636 69148
rect 345020 69096 345072 69148
rect 349804 69096 349856 69148
rect 356612 69096 356664 69148
rect 360844 69096 360896 69148
rect 104164 69028 104216 69080
rect 104900 69028 104952 69080
rect 117964 69028 118016 69080
rect 120540 69028 120592 69080
rect 162124 69028 162176 69080
rect 165252 69028 165304 69080
rect 210424 69028 210476 69080
rect 212540 69028 212592 69080
rect 224224 69028 224276 69080
rect 224960 69028 225012 69080
rect 229744 69028 229796 69080
rect 234804 69028 234856 69080
rect 242164 69028 242216 69080
rect 243912 69028 243964 69080
rect 269764 69028 269816 69080
rect 272064 69028 272116 69080
rect 279424 69028 279476 69080
rect 282000 69028 282052 69080
rect 288440 69028 288492 69080
rect 290280 69028 290332 69080
rect 298652 69028 298704 69080
rect 299756 69028 299808 69080
rect 300308 69028 300360 69080
rect 302240 69028 302292 69080
rect 304448 69028 304500 69080
rect 305644 69028 305696 69080
rect 307760 69028 307812 69080
rect 309784 69028 309836 69080
rect 312728 69028 312780 69080
rect 313924 69028 313976 69080
rect 316040 69028 316092 69080
rect 318064 69028 318116 69080
rect 330944 69028 330996 69080
rect 331864 69028 331916 69080
rect 348332 69028 348384 69080
rect 351184 69028 351236 69080
rect 355784 69028 355836 69080
rect 356704 69028 356756 69080
rect 357440 69028 357492 69080
rect 359464 69028 359516 69080
rect 362408 69028 362460 69080
rect 363604 69028 363656 69080
rect 366548 69028 366600 69080
rect 369124 69028 369176 69080
rect 398012 69028 398064 69080
rect 399484 69028 399536 69080
rect 438584 69028 438636 69080
rect 439504 69028 439556 69080
rect 443552 69028 443604 69080
rect 445024 69028 445076 69080
rect 455972 69028 456024 69080
rect 458824 69028 458876 69080
rect 460940 69028 460992 69080
rect 468484 69028 468536 69080
rect 470876 69028 470928 69080
rect 472624 69028 472676 69080
rect 475844 69028 475896 69080
rect 476764 69028 476816 69080
rect 480812 69028 480864 69080
rect 482284 69028 482336 69080
rect 207020 68416 207072 68468
rect 233240 68416 233292 68468
rect 253204 68416 253256 68468
rect 256332 68416 256384 68468
rect 149060 68348 149112 68400
rect 192576 68348 192628 68400
rect 193220 68348 193272 68400
rect 223212 68348 223264 68400
rect 370688 68348 370740 68400
rect 402980 68348 403032 68400
rect 434444 68348 434496 68400
rect 494152 68348 494204 68400
rect 7564 68280 7616 68332
rect 89076 68280 89128 68332
rect 93860 68280 93912 68332
rect 154580 68280 154632 68332
rect 171140 68280 171192 68332
rect 208400 68280 208452 68332
rect 227720 68280 227772 68332
rect 248052 68280 248104 68332
rect 249800 68280 249852 68332
rect 262956 68280 263008 68332
rect 383936 68280 383988 68332
rect 422300 68280 422352 68332
rect 465080 68280 465132 68332
rect 538220 68280 538272 68332
rect 489920 67600 489972 67652
rect 490196 67600 490248 67652
rect 209780 67056 209832 67108
rect 235632 67056 235684 67108
rect 200120 66988 200172 67040
rect 228180 66988 228232 67040
rect 80060 66920 80112 66972
rect 144552 66920 144604 66972
rect 165620 66920 165672 66972
rect 204260 66920 204312 66972
rect 4804 66852 4856 66904
rect 88340 66852 88392 66904
rect 115940 66852 115992 66904
rect 169392 66852 169444 66904
rect 175280 66852 175332 66904
rect 210792 66852 210844 66904
rect 238760 66852 238812 66904
rect 255504 66852 255556 66904
rect 375656 66852 375708 66904
rect 409880 66852 409932 66904
rect 479156 66852 479208 66904
rect 557540 66852 557592 66904
rect 255964 66240 256016 66292
rect 259644 66240 259696 66292
rect 324412 66172 324464 66224
rect 325056 66172 325108 66224
rect 224960 65764 225012 65816
rect 245660 65764 245712 65816
rect 196072 65628 196124 65680
rect 225696 65628 225748 65680
rect 259552 65628 259604 65680
rect 269580 65628 269632 65680
rect 44180 65492 44232 65544
rect 118884 65492 118936 65544
rect 157984 65492 158036 65544
rect 196716 65492 196768 65544
rect 211160 65492 211212 65544
rect 236460 65492 236512 65544
rect 245660 65492 245712 65544
rect 260472 65492 260524 65544
rect 402152 65492 402204 65544
rect 448520 65492 448572 65544
rect 484124 65492 484176 65544
rect 564532 65492 564584 65544
rect 146392 64336 146444 64388
rect 190460 64336 190512 64388
rect 220820 64336 220872 64388
rect 242992 64336 243044 64388
rect 84200 64200 84252 64252
rect 146484 64200 146536 64252
rect 192484 64200 192536 64252
rect 221004 64200 221056 64252
rect 29000 64132 29052 64184
rect 109040 64132 109092 64184
rect 189172 64132 189224 64184
rect 220912 64132 220964 64184
rect 242992 64132 243044 64184
rect 258080 64132 258132 64184
rect 481640 64132 481692 64184
rect 561680 64132 561732 64184
rect 121552 62908 121604 62960
rect 172612 62908 172664 62960
rect 444380 62840 444432 62892
rect 507860 62840 507912 62892
rect 46940 62772 46992 62824
rect 121644 62772 121696 62824
rect 178040 62772 178092 62824
rect 212632 62772 212684 62824
rect 214012 62772 214064 62824
rect 237472 62772 237524 62824
rect 478880 62772 478932 62824
rect 558920 62772 558972 62824
rect 484400 61344 484452 61396
rect 565820 61344 565872 61396
rect 577872 60664 577924 60716
rect 579988 60664 580040 60716
rect 13084 59984 13136 60036
rect 94228 59984 94280 60036
rect 3056 59304 3108 59356
rect 512092 59304 512144 59356
rect 74540 58692 74592 58744
rect 139492 58692 139544 58744
rect 27620 58624 27672 58676
rect 106648 58624 106700 58676
rect 174636 58624 174688 58676
rect 208584 58624 208636 58676
rect 469312 58624 469364 58676
rect 545120 58624 545172 58676
rect 67640 57264 67692 57316
rect 135352 57264 135404 57316
rect 429292 57264 429344 57316
rect 488632 57264 488684 57316
rect 17960 57196 18012 57248
rect 100760 57196 100812 57248
rect 182824 57196 182876 57248
rect 214104 57196 214156 57248
rect 473360 57196 473412 57248
rect 549260 57196 549312 57248
rect 30380 55836 30432 55888
rect 109224 55836 109276 55888
rect 144920 55836 144972 55888
rect 189448 55836 189500 55888
rect 415400 55836 415452 55888
rect 466552 55836 466604 55888
rect 487160 55836 487212 55888
rect 569960 55836 570012 55888
rect 433340 54544 433392 54596
rect 492680 54544 492732 54596
rect 44272 54476 44324 54528
rect 118700 54476 118752 54528
rect 490012 54476 490064 54528
rect 574100 54476 574152 54528
rect 41420 53048 41472 53100
rect 117320 53048 117372 53100
rect 491392 53048 491444 53100
rect 576124 53048 576176 53100
rect 37280 51688 37332 51740
rect 114652 51688 114704 51740
rect 151820 51688 151872 51740
rect 194600 51688 194652 51740
rect 440332 51688 440384 51740
rect 503720 51688 503772 51740
rect 102232 50396 102284 50448
rect 158812 50396 158864 50448
rect 24860 50328 24912 50380
rect 104992 50328 105044 50380
rect 188344 50328 188396 50380
rect 218152 50328 218204 50380
rect 439504 50328 439556 50380
rect 499580 50328 499632 50380
rect 92664 49036 92716 49088
rect 152188 49036 152240 49088
rect 425152 49036 425204 49088
rect 481640 49036 481692 49088
rect 49700 48968 49752 49020
rect 122932 48968 122984 49020
rect 218152 48968 218204 49020
rect 240140 48968 240192 49020
rect 449992 48968 450044 49020
rect 517520 48968 517572 49020
rect 512644 46860 512696 46912
rect 580172 46860 580224 46912
rect 60740 46180 60792 46232
rect 131212 46180 131264 46232
rect 400220 46180 400272 46232
rect 445760 46180 445812 46232
rect 445852 46180 445904 46232
rect 512092 46180 512144 46232
rect 110512 44888 110564 44940
rect 162124 44888 162176 44940
rect 431960 44888 432012 44940
rect 489920 44888 489972 44940
rect 53840 44820 53892 44872
rect 125692 44820 125744 44872
rect 223672 44820 223724 44872
rect 244280 44820 244332 44872
rect 379612 44820 379664 44872
rect 416872 44820 416924 44872
rect 458824 44820 458876 44872
rect 524420 44820 524472 44872
rect 63500 43460 63552 43512
rect 132500 43460 132552 43512
rect 436100 43460 436152 43512
rect 496820 43460 496872 43512
rect 17224 43392 17276 43444
rect 96712 43392 96764 43444
rect 142252 43392 142304 43444
rect 187700 43392 187752 43444
rect 476764 43392 476816 43444
rect 553400 43392 553452 43444
rect 56600 42100 56652 42152
rect 127072 42100 127124 42152
rect 8944 42032 8996 42084
rect 89812 42032 89864 42084
rect 102324 42032 102376 42084
rect 160192 42032 160244 42084
rect 231860 42032 231912 42084
rect 249892 42032 249944 42084
rect 419632 42032 419684 42084
rect 473360 42032 473412 42084
rect 481732 42032 481784 42084
rect 563060 42032 563112 42084
rect 99472 40740 99524 40792
rect 157340 40740 157392 40792
rect 52460 40672 52512 40724
rect 125600 40672 125652 40724
rect 436192 40672 436244 40724
rect 498200 40672 498252 40724
rect 111800 39448 111852 39500
rect 167000 39448 167052 39500
rect 423680 39380 423732 39432
rect 478880 39380 478932 39432
rect 34520 39312 34572 39364
rect 111892 39312 111944 39364
rect 477500 39312 477552 39364
rect 556252 39312 556304 39364
rect 85580 37952 85632 38004
rect 147772 37952 147824 38004
rect 432052 37952 432104 38004
rect 491392 37952 491444 38004
rect 35900 37884 35952 37936
rect 113272 37884 113324 37936
rect 485780 37884 485832 37936
rect 567200 37884 567252 37936
rect 26240 36524 26292 36576
rect 106372 36524 106424 36576
rect 118700 36524 118752 36576
rect 171324 36524 171376 36576
rect 445024 36524 445076 36576
rect 506480 36524 506532 36576
rect 98184 35164 98236 35216
rect 156052 35164 156104 35216
rect 430580 35164 430632 35216
rect 490012 35164 490064 35216
rect 31760 33736 31812 33788
rect 110604 33736 110656 33788
rect 114652 33736 114704 33788
rect 168380 33736 168432 33788
rect 427912 33736 427964 33788
rect 485780 33736 485832 33788
rect 490196 33736 490248 33788
rect 572720 33736 572772 33788
rect 3148 33056 3200 33108
rect 72424 33056 72476 33108
rect 514024 33056 514076 33108
rect 580172 33056 580224 33108
rect 417148 32444 417200 32496
rect 470692 32444 470744 32496
rect 107660 32376 107712 32428
rect 162952 32376 163004 32428
rect 453304 32376 453356 32428
rect 510620 32376 510672 32428
rect 91100 31016 91152 31068
rect 151912 31016 151964 31068
rect 156052 31016 156104 31068
rect 197544 31016 197596 31068
rect 390560 31016 390612 31068
rect 432052 31016 432104 31068
rect 454132 31016 454184 31068
rect 523040 31016 523092 31068
rect 60832 29588 60884 29640
rect 129832 29588 129884 29640
rect 135352 29588 135404 29640
rect 182180 29588 182232 29640
rect 412732 29588 412784 29640
rect 463792 29588 463844 29640
rect 471980 29588 472032 29640
rect 547880 29588 547932 29640
rect 86960 28228 87012 28280
rect 149152 28228 149204 28280
rect 151912 28228 151964 28280
rect 193588 28228 193640 28280
rect 382372 28228 382424 28280
rect 421012 28228 421064 28280
rect 425060 28228 425112 28280
rect 481732 28228 481784 28280
rect 73160 26868 73212 26920
rect 139400 26868 139452 26920
rect 147772 26868 147824 26920
rect 191932 26868 191984 26920
rect 409972 26868 410024 26920
rect 459652 26868 459704 26920
rect 466828 26868 466880 26920
rect 540980 26868 541032 26920
rect 134064 25576 134116 25628
rect 180892 25576 180944 25628
rect 69020 25508 69072 25560
rect 136640 25508 136692 25560
rect 367100 25508 367152 25560
rect 398840 25508 398892 25560
rect 407212 25508 407264 25560
rect 456892 25508 456944 25560
rect 462320 25508 462372 25560
rect 534080 25508 534132 25560
rect 55220 24080 55272 24132
rect 126980 24080 127032 24132
rect 127072 24080 127124 24132
rect 176752 24080 176804 24132
rect 404452 24080 404504 24132
rect 452752 24080 452804 24132
rect 456984 24080 457036 24132
rect 527180 24080 527232 24132
rect 420920 22788 420972 22840
rect 476212 22788 476264 22840
rect 40040 22720 40092 22772
rect 116032 22720 116084 22772
rect 129832 22720 129884 22772
rect 179420 22720 179472 22772
rect 365720 22720 365772 22772
rect 396264 22720 396316 22772
rect 456064 22720 456116 22772
rect 514760 22720 514812 22772
rect 175924 21428 175976 21480
rect 209872 21428 209924 21480
rect 22100 21360 22152 21412
rect 103520 21360 103572 21412
rect 103612 21360 103664 21412
rect 160100 21360 160152 21412
rect 161572 21360 161624 21412
rect 201592 21360 201644 21412
rect 378140 21360 378192 21412
rect 414112 21360 414164 21412
rect 419540 21360 419592 21412
rect 473544 21360 473596 21412
rect 474832 21360 474884 21412
rect 552020 21360 552072 21412
rect 3424 20612 3476 20664
rect 512000 20612 512052 20664
rect 577688 20612 577740 20664
rect 579804 20612 579856 20664
rect 157340 18640 157392 18692
rect 197452 18640 197504 18692
rect 372620 18640 372672 18692
rect 407212 18640 407264 18692
rect 100760 18572 100812 18624
rect 158720 18572 158772 18624
rect 392032 18572 392084 18624
rect 434812 18572 434864 18624
rect 451280 18572 451332 18624
rect 518900 18572 518952 18624
rect 399484 17348 399536 17400
rect 441712 17348 441764 17400
rect 162860 17280 162912 17332
rect 201500 17280 201552 17332
rect 57980 17212 58032 17264
rect 128360 17212 128412 17264
rect 143632 17212 143684 17264
rect 187884 17212 187936 17264
rect 383660 17212 383712 17264
rect 423680 17212 423732 17264
rect 441804 17212 441856 17264
rect 505100 17212 505152 17264
rect 158904 15988 158956 16040
rect 198832 15988 198884 16040
rect 139584 15920 139636 15972
rect 185308 15920 185360 15972
rect 427820 15920 427872 15972
rect 484768 15920 484820 15972
rect 51080 15852 51132 15904
rect 122840 15852 122892 15904
rect 123024 15852 123076 15904
rect 173900 15852 173952 15904
rect 329840 15852 329892 15904
rect 345296 15852 345348 15904
rect 353300 15852 353352 15904
rect 378416 15852 378468 15904
rect 389180 15852 389232 15904
rect 430856 15852 430908 15904
rect 459560 15852 459612 15904
rect 531320 15852 531372 15904
rect 386512 14560 386564 14612
rect 426808 14560 426860 14612
rect 422392 14492 422444 14544
rect 478144 14492 478196 14544
rect 69112 14424 69164 14476
rect 135260 14424 135312 14476
rect 135812 14424 135864 14476
rect 183560 14424 183612 14476
rect 183744 14424 183796 14476
rect 216680 14424 216732 14476
rect 345112 14424 345164 14476
rect 367744 14424 367796 14476
rect 394792 14424 394844 14476
rect 439136 14424 439188 14476
rect 476120 14424 476172 14476
rect 554780 14424 554832 14476
rect 351184 13336 351236 13388
rect 371332 13336 371384 13388
rect 371608 13200 371660 13252
rect 406016 13200 406068 13252
rect 150624 13132 150676 13184
rect 193312 13132 193364 13184
rect 387800 13132 387852 13184
rect 428464 13132 428516 13184
rect 132960 13064 133012 13116
rect 180800 13064 180852 13116
rect 205088 13064 205140 13116
rect 230572 13064 230624 13116
rect 360200 13064 360252 13116
rect 389456 13064 389508 13116
rect 403072 13064 403124 13116
rect 449808 13064 449860 13116
rect 470600 13064 470652 13116
rect 547972 13064 548024 13116
rect 345664 12996 345716 13048
rect 353576 12996 353628 13048
rect 338120 11840 338172 11892
rect 357532 11840 357584 11892
rect 137192 11772 137244 11824
rect 183836 11772 183888 11824
rect 342352 11772 342404 11824
rect 364616 11772 364668 11824
rect 367284 11772 367336 11824
rect 399024 11772 399076 11824
rect 24216 11704 24268 11756
rect 104164 11704 104216 11756
rect 128912 11704 128964 11756
rect 178132 11704 178184 11756
rect 186136 11704 186188 11756
rect 218060 11704 218112 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 259460 11704 259512 11756
rect 260656 11704 260708 11756
rect 356704 11704 356756 11756
rect 382372 11704 382424 11756
rect 391940 11704 391992 11756
rect 433984 11704 434036 11756
rect 438952 11704 439004 11756
rect 501328 11704 501380 11756
rect 363604 10412 363656 10464
rect 391112 10412 391164 10464
rect 111616 10344 111668 10396
rect 165712 10344 165764 10396
rect 178684 10344 178736 10396
rect 211252 10344 211304 10396
rect 332692 10344 332744 10396
rect 349160 10344 349212 10396
rect 364432 10344 364484 10396
rect 395344 10344 395396 10396
rect 429200 10344 429252 10396
rect 487160 10344 487212 10396
rect 65064 10276 65116 10328
rect 133880 10276 133932 10328
rect 164424 10276 164476 10328
rect 202880 10276 202932 10328
rect 342260 10276 342312 10328
rect 363512 10276 363564 10328
rect 378232 10276 378284 10328
rect 415492 10276 415544 10328
rect 473452 10276 473504 10328
rect 551008 10276 551060 10328
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 161296 9052 161348 9104
rect 200212 9052 200264 9104
rect 358820 9052 358872 9104
rect 388260 9052 388312 9104
rect 109316 8984 109368 9036
rect 164332 8984 164384 9036
rect 169576 8984 169628 9036
rect 206008 8984 206060 9036
rect 328460 8984 328512 9036
rect 343364 8984 343416 9036
rect 382280 8984 382332 9036
rect 420184 8984 420236 9036
rect 426440 8984 426492 9036
rect 484032 8984 484084 9036
rect 33600 8916 33652 8968
rect 110420 8916 110472 8968
rect 128176 8916 128228 8968
rect 176660 8916 176712 8968
rect 336832 8916 336884 8968
rect 356336 8916 356388 8968
rect 359464 8916 359516 8968
rect 384764 8916 384816 8968
rect 385132 8916 385184 8968
rect 424968 8916 425020 8968
rect 454040 8916 454092 8968
rect 523040 8916 523092 8968
rect 351920 7760 351972 7812
rect 377680 7760 377732 7812
rect 321652 7692 321704 7744
rect 335084 7692 335136 7744
rect 354680 7692 354732 7744
rect 381176 7692 381228 7744
rect 125876 7624 125928 7676
rect 175372 7624 175424 7676
rect 203892 7624 203944 7676
rect 230480 7624 230532 7676
rect 331864 7624 331916 7676
rect 346952 7624 347004 7676
rect 379520 7624 379572 7676
rect 416688 7624 416740 7676
rect 448612 7624 448664 7676
rect 515956 7624 516008 7676
rect 7656 7556 7708 7608
rect 92572 7556 92624 7608
rect 105728 7556 105780 7608
rect 161480 7556 161532 7608
rect 168380 7556 168432 7608
rect 205732 7556 205784 7608
rect 334348 7556 334400 7608
rect 352840 7556 352892 7608
rect 376852 7556 376904 7608
rect 413100 7556 413152 7608
rect 423864 7556 423916 7608
rect 480536 7556 480588 7608
rect 485872 7556 485924 7608
rect 569132 7556 569184 7608
rect 3424 6808 3476 6860
rect 511080 6808 511132 6860
rect 577504 6740 577556 6792
rect 579712 6740 579764 6792
rect 77392 6604 77444 6656
rect 142160 6604 142212 6656
rect 434720 6604 434772 6656
rect 495900 6604 495952 6656
rect 66720 6536 66772 6588
rect 134156 6536 134208 6588
rect 437480 6536 437532 6588
rect 499396 6536 499448 6588
rect 63224 6468 63276 6520
rect 131120 6468 131172 6520
rect 440240 6468 440292 6520
rect 502984 6468 503036 6520
rect 59636 6400 59688 6452
rect 129740 6400 129792 6452
rect 346492 6400 346544 6452
rect 370596 6400 370648 6452
rect 444472 6400 444524 6452
rect 510068 6400 510120 6452
rect 52552 6332 52604 6384
rect 124312 6332 124364 6384
rect 441620 6332 441672 6384
rect 506480 6332 506532 6384
rect 48964 6264 49016 6316
rect 121736 6264 121788 6316
rect 138848 6264 138900 6316
rect 185032 6264 185084 6316
rect 370044 6264 370096 6316
rect 402520 6264 402572 6316
rect 449900 6264 449952 6316
rect 517152 6264 517204 6316
rect 8760 6196 8812 6248
rect 93952 6196 94004 6248
rect 131764 6196 131816 6248
rect 179604 6196 179656 6248
rect 213368 6196 213420 6248
rect 237380 6196 237432 6248
rect 374184 6196 374236 6248
rect 409604 6196 409656 6248
rect 447140 6196 447192 6248
rect 513564 6196 513616 6248
rect 4068 6128 4120 6180
rect 89720 6128 89772 6180
rect 118792 6128 118844 6180
rect 171232 6128 171284 6180
rect 182548 6128 182600 6180
rect 215300 6128 215352 6180
rect 327080 6128 327132 6180
rect 342168 6128 342220 6180
rect 349252 6128 349304 6180
rect 374092 6128 374144 6180
rect 388168 6128 388220 6180
rect 429660 6128 429712 6180
rect 452660 6128 452712 6180
rect 520740 6128 520792 6180
rect 336096 5516 336148 5568
rect 339868 5516 339920 5568
rect 93952 5380 94004 5432
rect 153200 5380 153252 5432
rect 90364 5312 90416 5364
rect 150716 5312 150768 5364
rect 394700 5312 394752 5364
rect 437940 5312 437992 5364
rect 86868 5244 86920 5296
rect 147680 5244 147732 5296
rect 396172 5244 396224 5296
rect 441528 5244 441580 5296
rect 456800 5244 456852 5296
rect 526628 5244 526680 5296
rect 83280 5176 83332 5228
rect 146300 5176 146352 5228
rect 398932 5176 398984 5228
rect 445024 5176 445076 5228
rect 461032 5176 461084 5228
rect 533712 5176 533764 5228
rect 79692 5108 79744 5160
rect 143632 5108 143684 5160
rect 404360 5108 404412 5160
rect 452108 5108 452160 5160
rect 458180 5108 458232 5160
rect 530124 5108 530176 5160
rect 76196 5040 76248 5092
rect 140780 5040 140832 5092
rect 407120 5040 407172 5092
rect 455696 5040 455748 5092
rect 466460 5040 466512 5092
rect 540796 5040 540848 5092
rect 72608 4972 72660 5024
rect 138204 4972 138256 5024
rect 154212 4972 154264 5024
rect 195980 4972 196032 5024
rect 408868 4972 408920 5024
rect 459192 4972 459244 5024
rect 463700 4972 463752 5024
rect 537208 4972 537260 5024
rect 21824 4904 21876 4956
rect 102508 4904 102560 4956
rect 144736 4904 144788 4956
rect 189080 4904 189132 4956
rect 314660 4904 314712 4956
rect 324320 4904 324372 4956
rect 349804 4904 349856 4956
rect 367008 4904 367060 4956
rect 411352 4904 411404 4956
rect 462780 4904 462832 4956
rect 469220 4904 469272 4956
rect 544384 4904 544436 4956
rect 17040 4836 17092 4888
rect 99380 4836 99432 4888
rect 141240 4836 141292 4888
rect 186320 4836 186372 4888
rect 241704 4836 241756 4888
rect 256792 4836 256844 4888
rect 332600 4836 332652 4888
rect 349252 4836 349304 4888
rect 355324 4836 355376 4888
rect 375288 4836 375340 4888
rect 414020 4836 414072 4888
rect 466276 4836 466328 4888
rect 491300 4836 491352 4888
rect 576308 4836 576360 4888
rect 12348 4768 12400 4820
rect 96620 4768 96672 4820
rect 97448 4768 97500 4820
rect 155960 4768 156012 4820
rect 194416 4768 194468 4820
rect 223580 4768 223632 4820
rect 235816 4768 235868 4820
rect 252560 4768 252612 4820
rect 253480 4768 253532 4820
rect 265072 4768 265124 4820
rect 324412 4768 324464 4820
rect 338672 4768 338724 4820
rect 339592 4768 339644 4820
rect 359924 4768 359976 4820
rect 362960 4768 363012 4820
rect 393044 4768 393096 4820
rect 416780 4768 416832 4820
rect 469864 4768 469916 4820
rect 488540 4768 488592 4820
rect 572720 4768 572772 4820
rect 323584 4360 323636 4412
rect 328000 4360 328052 4412
rect 327724 4156 327776 4208
rect 331588 4156 331640 4208
rect 1676 4088 1728 4140
rect 7564 4088 7616 4140
rect 13544 4088 13596 4140
rect 17224 4088 17276 4140
rect 180248 4088 180300 4140
rect 182824 4088 182876 4140
rect 262956 4088 263008 4140
rect 269764 4088 269816 4140
rect 284300 4088 284352 4140
rect 287152 4088 287204 4140
rect 302332 4088 302384 4140
rect 303528 4088 303580 4140
rect 436744 4088 436796 4140
rect 443828 4088 443880 4140
rect 20628 4020 20680 4072
rect 28264 4020 28316 4072
rect 208584 4020 208636 4072
rect 221464 4020 221516 4072
rect 201500 3952 201552 4004
rect 217324 3952 217376 4004
rect 398104 3952 398156 4004
rect 408408 3952 408460 4004
rect 114008 3884 114060 3936
rect 156604 3884 156656 3936
rect 216864 3884 216916 3936
rect 235264 3884 235316 3936
rect 305644 3884 305696 3936
rect 309048 3884 309100 3936
rect 313924 3884 313976 3936
rect 320916 3884 320968 3936
rect 321560 3884 321612 3936
rect 333888 3884 333940 3936
rect 336004 3884 336056 3936
rect 351644 3884 351696 3936
rect 380900 3884 380952 3936
rect 418988 3884 419040 3936
rect 543004 3884 543056 3936
rect 557356 3884 557408 3936
rect 89168 3816 89220 3868
rect 140044 3816 140096 3868
rect 215668 3816 215720 3868
rect 233884 3816 233936 3868
rect 276020 3816 276072 3868
rect 278044 3816 278096 3868
rect 316132 3816 316184 3868
rect 326804 3816 326856 3868
rect 328552 3816 328604 3868
rect 344560 3816 344612 3868
rect 386420 3816 386472 3868
rect 426164 3816 426216 3868
rect 440884 3816 440936 3868
rect 450912 3816 450964 3868
rect 545764 3816 545816 3868
rect 564440 3816 564492 3868
rect 43076 3748 43128 3800
rect 50344 3748 50396 3800
rect 82084 3748 82136 3800
rect 135904 3748 135956 3800
rect 209872 3748 209924 3800
rect 229744 3748 229796 3800
rect 238116 3748 238168 3800
rect 247684 3748 247736 3800
rect 318892 3748 318944 3800
rect 330392 3748 330444 3800
rect 336740 3748 336792 3800
rect 355232 3748 355284 3800
rect 390652 3748 390704 3800
rect 433248 3748 433300 3800
rect 443644 3748 443696 3800
rect 458088 3748 458140 3800
rect 478236 3748 478288 3800
rect 539600 3748 539652 3800
rect 547144 3748 547196 3800
rect 571524 3748 571576 3800
rect 46664 3680 46716 3732
rect 117964 3680 118016 3732
rect 202696 3680 202748 3732
rect 225604 3680 225656 3732
rect 234620 3680 234672 3732
rect 246304 3680 246356 3732
rect 277124 3680 277176 3732
rect 279424 3680 279476 3732
rect 279516 3680 279568 3732
rect 283104 3680 283156 3732
rect 303712 3680 303764 3732
rect 307944 3680 307996 3732
rect 320272 3680 320324 3732
rect 332692 3680 332744 3732
rect 340880 3680 340932 3732
rect 361120 3680 361172 3732
rect 362224 3680 362276 3732
rect 372896 3680 372948 3732
rect 382924 3680 382976 3732
rect 391204 3680 391256 3732
rect 394240 3680 394292 3732
rect 396080 3680 396132 3732
rect 440332 3680 440384 3732
rect 446404 3680 446456 3732
rect 461584 3680 461636 3732
rect 468484 3680 468536 3732
rect 532516 3680 532568 3732
rect 548524 3680 548576 3732
rect 578608 3680 578660 3732
rect 39580 3612 39632 3664
rect 114560 3612 114612 3664
rect 195612 3612 195664 3664
rect 224224 3612 224276 3664
rect 231032 3612 231084 3664
rect 242256 3612 242308 3664
rect 305000 3612 305052 3664
rect 310244 3612 310296 3664
rect 313648 3612 313700 3664
rect 323308 3612 323360 3664
rect 324596 3612 324648 3664
rect 337476 3612 337528 3664
rect 338488 3612 338540 3664
rect 358728 3612 358780 3664
rect 360844 3612 360896 3664
rect 383568 3612 383620 3664
rect 390652 3612 390704 3664
rect 400588 3612 400640 3664
rect 447416 3612 447468 3664
rect 450544 3612 450596 3664
rect 468668 3612 468720 3664
rect 472624 3612 472676 3664
rect 546684 3612 546736 3664
rect 549904 3612 549956 3664
rect 582196 3612 582248 3664
rect 5264 3476 5316 3528
rect 10324 3544 10376 3596
rect 15936 3544 15988 3596
rect 98092 3544 98144 3596
rect 117596 3544 117648 3596
rect 164884 3544 164936 3596
rect 181444 3544 181496 3596
rect 9956 3476 10008 3528
rect 13084 3476 13136 3528
rect 14740 3476 14792 3528
rect 98000 3476 98052 3528
rect 118700 3476 118752 3528
rect 119896 3476 119948 3528
rect 121092 3476 121144 3528
rect 167644 3476 167696 3528
rect 173164 3476 173216 3528
rect 174636 3476 174688 3528
rect 176660 3476 176712 3528
rect 178684 3476 178736 3528
rect 187332 3476 187384 3528
rect 188344 3476 188396 3528
rect 188528 3544 188580 3596
rect 219532 3544 219584 3596
rect 227536 3544 227588 3596
rect 239404 3544 239456 3596
rect 251180 3544 251232 3596
rect 252376 3544 252428 3596
rect 258264 3544 258316 3596
rect 261484 3544 261536 3596
rect 267740 3544 267792 3596
rect 268476 3544 268528 3596
rect 283104 3544 283156 3596
rect 285772 3544 285824 3596
rect 317788 3544 317840 3596
rect 329196 3544 329248 3596
rect 331312 3544 331364 3596
rect 348056 3544 348108 3596
rect 350908 3544 350960 3596
rect 376484 3544 376536 3596
rect 377404 3544 377456 3596
rect 387156 3544 387208 3596
rect 405740 3544 405792 3596
rect 454500 3544 454552 3596
rect 482284 3544 482336 3596
rect 560852 3544 560904 3596
rect 213920 3476 213972 3528
rect 226340 3476 226392 3528
rect 228364 3476 228416 3528
rect 6460 3408 6512 3460
rect 92480 3408 92532 3460
rect 96252 3408 96304 3460
rect 144184 3408 144236 3460
rect 160100 3408 160152 3460
rect 28908 3340 28960 3392
rect 32404 3340 32456 3392
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 69020 3340 69072 3392
rect 69940 3340 69992 3392
rect 174268 3408 174320 3460
rect 175924 3408 175976 3460
rect 177856 3408 177908 3460
rect 210424 3408 210476 3460
rect 219256 3408 219308 3460
rect 174544 3340 174596 3392
rect 190828 3340 190880 3392
rect 192484 3340 192536 3392
rect 209780 3340 209832 3392
rect 210976 3340 211028 3392
rect 2872 3272 2924 3324
rect 8944 3272 8996 3324
rect 19432 3272 19484 3324
rect 25504 3272 25556 3324
rect 222752 3340 222804 3392
rect 242164 3476 242216 3528
rect 245200 3476 245252 3528
rect 255964 3476 256016 3528
rect 272432 3476 272484 3528
rect 273904 3476 273956 3528
rect 300952 3476 301004 3528
rect 305552 3476 305604 3528
rect 309784 3476 309836 3528
rect 313832 3476 313884 3528
rect 323032 3476 323084 3528
rect 336280 3476 336332 3528
rect 341064 3476 341116 3528
rect 362316 3476 362368 3528
rect 369124 3476 369176 3528
rect 397736 3476 397788 3528
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 400864 3476 400916 3528
rect 411904 3476 411956 3528
rect 412640 3476 412692 3528
rect 465172 3476 465224 3528
rect 473360 3476 473412 3528
rect 474188 3476 474240 3528
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 494060 3476 494112 3528
rect 581000 3476 581052 3528
rect 238024 3408 238076 3460
rect 240508 3408 240560 3460
rect 253204 3408 253256 3460
rect 290188 3408 290240 3460
rect 291200 3408 291252 3460
rect 296812 3408 296864 3460
rect 299664 3408 299716 3460
rect 307024 3408 307076 3460
rect 311440 3408 311492 3460
rect 313372 3408 313424 3460
rect 322112 3408 322164 3460
rect 326068 3408 326120 3460
rect 340972 3408 341024 3460
rect 349160 3408 349212 3460
rect 350448 3408 350500 3460
rect 310520 3340 310572 3392
rect 318524 3340 318576 3392
rect 346584 3340 346636 3392
rect 369400 3408 369452 3460
rect 371240 3408 371292 3460
rect 404820 3408 404872 3460
rect 418252 3408 418304 3460
rect 472256 3408 472308 3460
rect 495532 3408 495584 3460
rect 583392 3408 583444 3460
rect 435364 3340 435416 3392
rect 436744 3340 436796 3392
rect 547880 3340 547932 3392
rect 548708 3340 548760 3392
rect 311164 3272 311216 3324
rect 315028 3272 315080 3324
rect 318064 3272 318116 3324
rect 325608 3272 325660 3324
rect 358084 3272 358136 3324
rect 365812 3272 365864 3324
rect 374644 3272 374696 3324
rect 379980 3272 380032 3324
rect 11152 3204 11204 3256
rect 14464 3204 14516 3256
rect 309324 3204 309376 3256
rect 316224 3204 316276 3256
rect 576124 3204 576176 3256
rect 577412 3204 577464 3256
rect 35992 3136 36044 3188
rect 39304 3136 39356 3188
rect 167184 3136 167236 3188
rect 170404 3136 170456 3188
rect 540244 3136 540296 3188
rect 543188 3136 543240 3188
rect 572 3068 624 3120
rect 4804 3068 4856 3120
rect 309140 3068 309192 3120
rect 317328 3068 317380 3120
rect 155408 3000 155460 3052
rect 157984 3000 158036 3052
rect 295432 3000 295484 3052
rect 297272 3000 297324 3052
rect 303528 3000 303580 3052
rect 306748 3000 306800 3052
rect 296904 2932 296956 2984
rect 298468 2932 298520 2984
rect 306472 2932 306524 2984
rect 312636 2932 312688 2984
rect 393964 2932 394016 2984
rect 401324 2932 401376 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 7564 637832 7616 637838
rect 7564 637774 7616 637780
rect 3516 634908 3568 634914
rect 3516 634850 3568 634856
rect 3424 633616 3476 633622
rect 3424 633558 3476 633564
rect 3332 632596 3384 632602
rect 3332 632538 3384 632544
rect 3240 632392 3292 632398
rect 3240 632334 3292 632340
rect 3148 619608 3200 619614
rect 3148 619550 3200 619556
rect 3160 619177 3188 619550
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 2780 607096 2832 607102
rect 2780 607038 2832 607044
rect 2792 606121 2820 607038
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 3148 580984 3200 580990
rect 3148 580926 3200 580932
rect 3160 580009 3188 580926
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3252 566953 3280 632334
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3344 553897 3372 632538
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3332 528556 3384 528562
rect 3332 528498 3384 528504
rect 3344 527921 3372 528498
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3332 501832 3384 501838
rect 3330 501800 3332 501809
rect 3384 501800 3386 501809
rect 3330 501735 3386 501744
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3344 475697 3372 476002
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3332 463684 3384 463690
rect 3332 463626 3384 463632
rect 3344 462641 3372 463626
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 2780 372360 2832 372366
rect 2780 372302 2832 372308
rect 2792 371385 2820 372302
rect 2778 371376 2834 371385
rect 2778 371311 2834 371320
rect 2964 346384 3016 346390
rect 2964 346326 3016 346332
rect 2976 345409 3004 346326
rect 2962 345400 3018 345409
rect 2962 345335 3018 345344
rect 2780 319864 2832 319870
rect 2780 319806 2832 319812
rect 2792 319297 2820 319806
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 2780 254992 2832 254998
rect 2780 254934 2832 254940
rect 2792 254153 2820 254934
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3436 188873 3464 633558
rect 3528 632097 3556 634850
rect 4068 633888 4120 633894
rect 4068 633830 4120 633836
rect 3884 633820 3936 633826
rect 3884 633762 3936 633768
rect 3792 633752 3844 633758
rect 3792 633694 3844 633700
rect 3700 632800 3752 632806
rect 3700 632742 3752 632748
rect 3608 632188 3660 632194
rect 3608 632130 3660 632136
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 631272 3570 631281
rect 3514 631207 3570 631216
rect 3528 201929 3556 631207
rect 3620 241097 3648 632130
rect 3712 293185 3740 632742
rect 3804 306241 3832 633694
rect 3896 358465 3924 633762
rect 3976 632256 4028 632262
rect 3976 632198 4028 632204
rect 3988 449585 4016 632198
rect 4080 514865 4108 633830
rect 4988 633684 5040 633690
rect 4988 633626 5040 633632
rect 4896 633548 4948 633554
rect 4896 633490 4948 633496
rect 4804 633480 4856 633486
rect 4804 633422 4856 633428
rect 4066 514856 4122 514865
rect 4066 514791 4122 514800
rect 3974 449576 4030 449585
rect 3974 449511 4030 449520
rect 3882 358456 3938 358465
rect 3882 358391 3938 358400
rect 3790 306232 3846 306241
rect 3790 306167 3846 306176
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3606 241088 3662 241097
rect 3606 241023 3662 241032
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 2780 149932 2832 149938
rect 2780 149874 2832 149880
rect 2792 149841 2820 149874
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4816 97782 4844 633422
rect 4908 149938 4936 633490
rect 5000 254998 5028 633626
rect 5264 632936 5316 632942
rect 5264 632878 5316 632884
rect 5172 630828 5224 630834
rect 5172 630770 5224 630776
rect 5080 630760 5132 630766
rect 5080 630702 5132 630708
rect 5092 319870 5120 630702
rect 5184 372366 5212 630770
rect 5276 607102 5304 632878
rect 5264 607096 5316 607102
rect 5264 607038 5316 607044
rect 7576 501838 7604 637774
rect 13084 637764 13136 637770
rect 13084 637706 13136 637712
rect 7564 501832 7616 501838
rect 7564 501774 7616 501780
rect 13096 398818 13124 637706
rect 40052 637090 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 71792 638450 71820 702986
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 105464 696250 105492 703520
rect 137848 697610 137876 703520
rect 154132 700670 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 137836 697604 137888 697610
rect 137836 697546 137888 697552
rect 105452 696244 105504 696250
rect 105452 696186 105504 696192
rect 71780 638444 71832 638450
rect 71780 638386 71832 638392
rect 68376 638308 68428 638314
rect 68376 638250 68428 638256
rect 58624 638172 58676 638178
rect 58624 638114 58676 638120
rect 57244 637968 57296 637974
rect 57244 637910 57296 637916
rect 40040 637084 40092 637090
rect 40040 637026 40092 637032
rect 53104 636880 53156 636886
rect 53104 636822 53156 636828
rect 21364 636336 21416 636342
rect 21364 636278 21416 636284
rect 13084 398812 13136 398818
rect 13084 398754 13136 398760
rect 5172 372360 5224 372366
rect 5172 372302 5224 372308
rect 5080 319864 5132 319870
rect 5080 319806 5132 319812
rect 4988 254992 5040 254998
rect 4988 254934 5040 254940
rect 21376 215286 21404 636278
rect 53116 411262 53144 636822
rect 53104 411256 53156 411262
rect 53104 411198 53156 411204
rect 57256 346390 57284 637910
rect 58636 463690 58664 638114
rect 66904 636744 66956 636750
rect 66904 636686 66956 636692
rect 64144 636540 64196 636546
rect 64144 636482 64196 636488
rect 62764 635044 62816 635050
rect 62764 634986 62816 634992
rect 62776 476066 62804 634986
rect 62764 476060 62816 476066
rect 62764 476002 62816 476008
rect 58624 463684 58676 463690
rect 58624 463626 58676 463632
rect 57244 346384 57296 346390
rect 57244 346326 57296 346332
rect 21364 215280 21416 215286
rect 21364 215222 21416 215228
rect 4896 149932 4948 149938
rect 4896 149874 4948 149880
rect 64156 111790 64184 636482
rect 66916 267714 66944 636686
rect 68284 636472 68336 636478
rect 68284 636414 68336 636420
rect 66904 267708 66956 267714
rect 66904 267650 66956 267656
rect 64144 111784 64196 111790
rect 64144 111726 64196 111732
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 68296 71738 68324 636414
rect 68388 619614 68416 638250
rect 161848 638036 161900 638042
rect 161848 637978 161900 637984
rect 150532 637900 150584 637906
rect 150532 637842 150584 637848
rect 109040 637696 109092 637702
rect 109040 637638 109092 637644
rect 105268 637628 105320 637634
rect 105268 637570 105320 637576
rect 71044 636608 71096 636614
rect 71044 636550 71096 636556
rect 68376 619608 68428 619614
rect 68376 619550 68428 619556
rect 71056 164218 71084 636550
rect 72424 636404 72476 636410
rect 72424 636346 72476 636352
rect 71320 635316 71372 635322
rect 71320 635258 71372 635264
rect 71228 635180 71280 635186
rect 71228 635122 71280 635128
rect 71136 634976 71188 634982
rect 71136 634918 71188 634924
rect 71148 423638 71176 634918
rect 71240 528562 71268 635122
rect 71332 580990 71360 635258
rect 71320 580984 71372 580990
rect 71320 580926 71372 580932
rect 71228 528556 71280 528562
rect 71228 528498 71280 528504
rect 71136 423632 71188 423638
rect 71136 423574 71188 423580
rect 71044 164212 71096 164218
rect 71044 164154 71096 164160
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 68284 71732 68336 71738
rect 68284 71674 68336 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 50344 70168 50396 70174
rect 50344 70110 50396 70116
rect 39304 70032 39356 70038
rect 39304 69974 39356 69980
rect 28264 69964 28316 69970
rect 28264 69906 28316 69912
rect 25504 69828 25556 69834
rect 25504 69770 25556 69776
rect 14464 69760 14516 69766
rect 14464 69702 14516 69708
rect 10324 69692 10376 69698
rect 10324 69634 10376 69640
rect 7564 68332 7616 68338
rect 7564 68274 7616 68280
rect 4804 66904 4856 66910
rect 4804 66846 4856 66852
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 584 480 612 3062
rect 1688 480 1716 4082
rect 2872 3324 2924 3330
rect 2872 3266 2924 3272
rect 2884 480 2912 3266
rect 4080 480 4108 6122
rect 4816 3126 4844 66846
rect 7576 4146 7604 68274
rect 8944 42084 8996 42090
rect 8944 42026 8996 42032
rect 7656 7608 7708 7614
rect 7656 7550 7708 7556
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 5276 480 5304 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 7550
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8772 480 8800 6190
rect 8956 3330 8984 42026
rect 10336 3602 10364 69634
rect 13084 60036 13136 60042
rect 13084 59978 13136 59984
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 8944 3324 8996 3330
rect 8944 3266 8996 3272
rect 9968 480 9996 3470
rect 11152 3256 11204 3262
rect 11152 3198 11204 3204
rect 11164 480 11192 3198
rect 12360 480 12388 4762
rect 13096 3534 13124 59978
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13556 480 13584 4082
rect 14476 3262 14504 69702
rect 17960 57248 18012 57254
rect 17960 57190 18012 57196
rect 17224 43444 17276 43450
rect 17224 43386 17276 43392
rect 17040 4888 17092 4894
rect 17040 4830 17092 4836
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14464 3256 14516 3262
rect 14464 3198 14516 3204
rect 14752 480 14780 3470
rect 15948 480 15976 3538
rect 17052 480 17080 4830
rect 17236 4146 17264 43386
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 57190
rect 24860 50380 24912 50386
rect 24860 50322 24912 50328
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22112 16574 22140 21354
rect 24872 16574 24900 50322
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 21824 4956 21876 4962
rect 21824 4898 21876 4904
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 19432 3324 19484 3330
rect 19432 3266 19484 3272
rect 19444 480 19472 3266
rect 20640 480 20668 4014
rect 21836 480 21864 4898
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24228 480 24256 11698
rect 25332 480 25360 16546
rect 25516 3330 25544 69770
rect 27620 58676 27672 58682
rect 27620 58618 27672 58624
rect 26240 36576 26292 36582
rect 26240 36518 26292 36524
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 36518
rect 27632 16574 27660 58618
rect 27632 16546 27752 16574
rect 27724 480 27752 16546
rect 28276 4078 28304 69906
rect 32404 69896 32456 69902
rect 32404 69838 32456 69844
rect 29000 64184 29052 64190
rect 29000 64126 29052 64132
rect 29012 16574 29040 64126
rect 30380 55888 30432 55894
rect 30380 55830 30432 55836
rect 30392 16574 30420 55830
rect 31760 33788 31812 33794
rect 31760 33730 31812 33736
rect 31772 16574 31800 33730
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3398 32444 69838
rect 37280 51740 37332 51746
rect 37280 51682 37332 51688
rect 34520 39364 34572 39370
rect 34520 39306 34572 39312
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33612 480 33640 8910
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 39306
rect 35900 37936 35952 37942
rect 35900 37878 35952 37884
rect 35912 16574 35940 37878
rect 37292 16574 37320 51682
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 36004 480 36032 3130
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 39316 3194 39344 69974
rect 44180 65544 44232 65550
rect 44180 65486 44232 65492
rect 41420 53100 41472 53106
rect 41420 53042 41472 53048
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40052 16574 40080 22714
rect 41432 16574 41460 53042
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39592 480 39620 3606
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 44192 6914 44220 65486
rect 46940 62824 46992 62830
rect 46940 62766 46992 62772
rect 44272 54528 44324 54534
rect 44272 54470 44324 54476
rect 44284 16574 44312 54470
rect 46952 16574 46980 62766
rect 49700 49020 49752 49026
rect 49700 48962 49752 48968
rect 49712 16574 49740 48962
rect 44284 16546 45048 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 43088 480 43116 3742
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 46676 480 46704 3674
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 6316 49016 6322
rect 48964 6258 49016 6264
rect 48976 480 49004 6258
rect 50172 480 50200 16546
rect 50356 3806 50384 70110
rect 70400 70100 70452 70106
rect 70400 70042 70452 70048
rect 67640 57316 67692 57322
rect 67640 57258 67692 57264
rect 60740 46232 60792 46238
rect 60740 46174 60792 46180
rect 53840 44872 53892 44878
rect 53840 44814 53892 44820
rect 52460 40724 52512 40730
rect 52460 40666 52512 40672
rect 52472 16574 52500 40666
rect 53852 16574 53880 44814
rect 56600 42152 56652 42158
rect 56600 42094 56652 42100
rect 55220 24132 55272 24138
rect 55220 24074 55272 24080
rect 55232 16574 55260 24074
rect 56612 16574 56640 42094
rect 57980 17264 58032 17270
rect 57980 17206 58032 17212
rect 57992 16574 58020 17206
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 51080 15904 51132 15910
rect 51080 15846 51132 15852
rect 50344 3800 50396 3806
rect 50344 3742 50396 3748
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 15846
rect 52552 6384 52604 6390
rect 52552 6326 52604 6332
rect 52564 480 52592 6326
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 59636 6452 59688 6458
rect 59636 6394 59688 6400
rect 59648 480 59676 6394
rect 60752 3398 60780 46174
rect 63500 43512 63552 43518
rect 63500 43454 63552 43460
rect 60832 29640 60884 29646
rect 60832 29582 60884 29588
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 29582
rect 63512 16574 63540 43454
rect 63512 16546 64368 16574
rect 63224 6520 63276 6526
rect 63224 6462 63276 6468
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 6462
rect 64340 480 64368 16546
rect 65064 10328 65116 10334
rect 65064 10270 65116 10276
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 10270
rect 66720 6588 66772 6594
rect 66720 6530 66772 6536
rect 66732 480 66760 6530
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 57258
rect 69020 25560 69072 25566
rect 69020 25502 69072 25508
rect 69032 3398 69060 25502
rect 70412 16574 70440 70042
rect 72436 33114 72464 636346
rect 82726 636304 82782 636313
rect 82726 636239 82782 636248
rect 94228 636268 94280 636274
rect 79138 633448 79194 633457
rect 79138 633383 79194 633392
rect 79152 631938 79180 633383
rect 82740 631938 82768 636239
rect 94228 636210 94280 636216
rect 90454 634944 90510 634953
rect 90454 634879 90510 634888
rect 86682 633584 86738 633593
rect 86682 633519 86738 633528
rect 86696 631938 86724 633519
rect 90468 631938 90496 634879
rect 94240 631938 94268 636210
rect 97906 633856 97962 633865
rect 97906 633791 97962 633800
rect 97920 631938 97948 633791
rect 105280 631938 105308 637570
rect 109052 631938 109080 637638
rect 147036 636812 147088 636818
rect 147036 636754 147088 636760
rect 124128 636676 124180 636682
rect 124128 636618 124180 636624
rect 113088 634840 113140 634846
rect 113088 634782 113140 634788
rect 113100 631938 113128 634782
rect 120630 632360 120686 632369
rect 120630 632295 120686 632304
rect 116858 632088 116914 632097
rect 116858 632023 116914 632032
rect 116872 631938 116900 632023
rect 120644 631938 120672 632295
rect 124140 631938 124168 636618
rect 139308 634296 139360 634302
rect 139308 634238 139360 634244
rect 131948 633956 132000 633962
rect 131948 633898 132000 633904
rect 127854 632120 127906 632126
rect 127854 632062 127906 632068
rect 78844 631910 79180 631938
rect 82616 631910 82768 631938
rect 86388 631910 86724 631938
rect 90160 631910 90496 631938
rect 93932 631910 94268 631938
rect 97704 631910 97948 631938
rect 105248 631910 105308 631938
rect 109020 631910 109080 631938
rect 112792 631910 113128 631938
rect 116564 631910 116900 631938
rect 120336 631910 120672 631938
rect 124108 631910 124168 631938
rect 127866 631924 127894 632062
rect 131960 631938 131988 633898
rect 135720 632460 135772 632466
rect 135720 632402 135772 632408
rect 135732 631938 135760 632402
rect 139320 631938 139348 634238
rect 147048 631938 147076 636754
rect 150544 631938 150572 637842
rect 154488 634024 154540 634030
rect 154488 633966 154540 633972
rect 154500 631938 154528 633966
rect 158352 632868 158404 632874
rect 158352 632810 158404 632816
rect 158364 631938 158392 632810
rect 161860 631938 161888 637978
rect 169772 637158 169800 702406
rect 201512 642394 201540 702986
rect 218992 700806 219020 703520
rect 218980 700800 219032 700806
rect 218980 700742 219032 700748
rect 229744 643136 229796 643142
rect 229744 643078 229796 643084
rect 201500 642388 201552 642394
rect 201500 642330 201552 642336
rect 184480 638240 184532 638246
rect 184480 638182 184532 638188
rect 173164 638104 173216 638110
rect 173164 638046 173216 638052
rect 169760 637152 169812 637158
rect 169760 637094 169812 637100
rect 165896 634092 165948 634098
rect 165896 634034 165948 634040
rect 165908 631938 165936 634034
rect 173176 631938 173204 638046
rect 180708 636948 180760 636954
rect 180708 636890 180760 636896
rect 177212 634228 177264 634234
rect 177212 634170 177264 634176
rect 177224 631938 177252 634170
rect 180720 631938 180748 636890
rect 184492 631938 184520 638182
rect 226248 635452 226300 635458
rect 226248 635394 226300 635400
rect 214932 635384 214984 635390
rect 214932 635326 214984 635332
rect 203616 635248 203668 635254
rect 203616 635190 203668 635196
rect 199844 635112 199896 635118
rect 199844 635054 199896 635060
rect 192300 634160 192352 634166
rect 192300 634102 192352 634108
rect 192312 631938 192340 634102
rect 195888 632324 195940 632330
rect 195888 632266 195940 632272
rect 195900 631938 195928 632266
rect 199856 631938 199884 635054
rect 203628 631938 203656 635190
rect 207388 632528 207440 632534
rect 207388 632470 207440 632476
rect 207400 631938 207428 632470
rect 214944 631938 214972 635326
rect 216680 634364 216732 634370
rect 216680 634306 216732 634312
rect 216692 632806 216720 634306
rect 216680 632800 216732 632806
rect 216680 632742 216732 632748
rect 222476 632800 222528 632806
rect 222476 632742 222528 632748
rect 218704 632664 218756 632670
rect 218704 632606 218756 632612
rect 218716 631938 218744 632606
rect 222488 631938 222516 632742
rect 226260 631938 226288 635394
rect 229756 631938 229784 643078
rect 234632 641034 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267464 700596 267516 700602
rect 267464 700538 267516 700544
rect 256148 700460 256200 700466
rect 256148 700402 256200 700408
rect 241060 696992 241112 696998
rect 241060 696934 241112 696940
rect 237288 670812 237340 670818
rect 237288 670754 237340 670760
rect 234620 641028 234672 641034
rect 234620 640970 234672 640976
rect 237300 631938 237328 670754
rect 241072 631938 241100 696934
rect 244832 683256 244884 683262
rect 244832 683198 244884 683204
rect 244844 631938 244872 683198
rect 252376 638376 252428 638382
rect 252376 638318 252428 638324
rect 248880 637016 248932 637022
rect 248880 636958 248932 636964
rect 248892 631938 248920 636958
rect 252388 631938 252416 638318
rect 256160 631938 256188 700402
rect 263692 639600 263744 639606
rect 263692 639542 263744 639548
rect 260196 635520 260248 635526
rect 260196 635462 260248 635468
rect 260208 631938 260236 635462
rect 263704 631938 263732 639542
rect 267476 631938 267504 700538
rect 267660 699038 267688 703520
rect 283852 700942 283880 703520
rect 283840 700936 283892 700942
rect 283840 700878 283892 700884
rect 290096 700868 290148 700874
rect 290096 700810 290148 700816
rect 278780 700732 278832 700738
rect 278780 700674 278832 700680
rect 267648 699032 267700 699038
rect 267648 698974 267700 698980
rect 275008 698964 275060 698970
rect 275008 698906 275060 698912
rect 271512 635588 271564 635594
rect 271512 635530 271564 635536
rect 271524 631938 271552 635530
rect 275020 631938 275048 698906
rect 278792 631938 278820 700674
rect 286324 663060 286376 663066
rect 286324 663002 286376 663008
rect 282828 635656 282880 635662
rect 282828 635598 282880 635604
rect 282840 631938 282868 635598
rect 286336 631938 286364 663002
rect 290108 631938 290136 700810
rect 297640 699032 297692 699038
rect 297640 698974 297692 698980
rect 293868 635724 293920 635730
rect 293868 635666 293920 635672
rect 293880 631938 293908 635666
rect 297652 631938 297680 698974
rect 299492 635730 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 301412 700936 301464 700942
rect 301412 700878 301464 700884
rect 299480 635724 299532 635730
rect 299480 635666 299532 635672
rect 301424 631938 301452 700878
rect 312728 700800 312780 700806
rect 312728 700742 312780 700748
rect 308956 642388 309008 642394
rect 308956 642330 309008 642336
rect 305184 641028 305236 641034
rect 305184 640970 305236 640976
rect 305196 631938 305224 640970
rect 308968 631938 308996 642330
rect 312740 631938 312768 700742
rect 324044 700664 324096 700670
rect 324044 700606 324096 700612
rect 320272 697604 320324 697610
rect 320272 697546 320324 697552
rect 316132 637152 316184 637158
rect 316132 637094 316184 637100
rect 131652 631910 131988 631938
rect 135424 631910 135760 631938
rect 139196 631910 139348 631938
rect 146740 631910 147076 631938
rect 150512 631910 150572 631938
rect 154284 631910 154528 631938
rect 158056 631910 158392 631938
rect 161828 631910 161888 631938
rect 165600 631910 165936 631938
rect 173144 631910 173204 631938
rect 176916 631910 177252 631938
rect 180688 631910 180748 631938
rect 184460 631910 184520 631938
rect 192004 631910 192340 631938
rect 195776 631910 195928 631938
rect 199548 631910 199884 631938
rect 203320 631910 203656 631938
rect 207092 631910 207428 631938
rect 214636 631910 214972 631938
rect 218408 631910 218744 631938
rect 222180 631910 222516 631938
rect 225952 631910 226288 631938
rect 229724 631910 229784 631938
rect 237268 631910 237328 631938
rect 241040 631910 241100 631938
rect 244812 631910 244872 631938
rect 248584 631910 248920 631938
rect 252356 631910 252416 631938
rect 256128 631910 256188 631938
rect 259900 631910 260236 631938
rect 263672 631910 263732 631938
rect 267444 631910 267504 631938
rect 271216 631910 271552 631938
rect 274988 631910 275048 631938
rect 278760 631910 278820 631938
rect 282532 631910 282868 631938
rect 286304 631910 286364 631938
rect 290076 631910 290136 631938
rect 293848 631910 293908 631938
rect 297620 631910 297680 631938
rect 301392 631910 301452 631938
rect 305164 631910 305224 631938
rect 308936 631910 308996 631938
rect 312708 631910 312768 631938
rect 316144 631938 316172 637094
rect 320284 631938 320312 697546
rect 324056 631938 324084 700606
rect 327816 696244 327868 696250
rect 327816 696186 327868 696192
rect 327828 631938 327856 696186
rect 331232 663066 331260 702986
rect 348804 700874 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700868 348844 700874
rect 348792 700810 348844 700816
rect 335360 700528 335412 700534
rect 335360 700470 335412 700476
rect 331220 663060 331272 663066
rect 331220 663002 331272 663008
rect 331588 638444 331640 638450
rect 331588 638386 331640 638392
rect 331600 631938 331628 638386
rect 335372 631938 335400 700470
rect 346676 700392 346728 700398
rect 346676 700334 346728 700340
rect 342904 700324 342956 700330
rect 342904 700266 342956 700272
rect 338764 637084 338816 637090
rect 338764 637026 338816 637032
rect 316144 631910 316480 631938
rect 320252 631910 320312 631938
rect 324024 631910 324084 631938
rect 327796 631910 327856 631938
rect 331568 631910 331628 631938
rect 335340 631910 335400 631938
rect 338776 631938 338804 637026
rect 342916 631938 342944 700266
rect 346688 631938 346716 700334
rect 350448 683188 350500 683194
rect 350448 683130 350500 683136
rect 350460 631938 350488 683130
rect 357992 670744 358044 670750
rect 357992 670686 358044 670692
rect 354220 656940 354272 656946
rect 354220 656882 354272 656888
rect 354232 631938 354260 656882
rect 358004 631938 358032 670686
rect 364352 635662 364380 702406
rect 397472 698970 397500 703520
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 397460 698964 397512 698970
rect 397460 698906 397512 698912
rect 369308 638308 369360 638314
rect 369308 638250 369360 638256
rect 364340 635656 364392 635662
rect 364340 635598 364392 635604
rect 361580 634908 361632 634914
rect 361580 634850 361632 634856
rect 338776 631910 339112 631938
rect 342884 631910 342944 631938
rect 346656 631910 346716 631938
rect 350428 631910 350488 631938
rect 354200 631910 354260 631938
rect 357972 631910 358032 631938
rect 361592 631938 361620 634850
rect 365628 634296 365680 634302
rect 365628 634238 365680 634244
rect 366548 634296 366600 634302
rect 366548 634238 366600 634244
rect 365168 632936 365220 632942
rect 365168 632878 365220 632884
rect 365180 631938 365208 632878
rect 365640 632738 365668 634238
rect 365628 632732 365680 632738
rect 365628 632674 365680 632680
rect 361592 631910 361744 631938
rect 365180 631910 365516 631938
rect 142804 631576 142856 631582
rect 142804 631518 142856 631524
rect 146944 631576 146996 631582
rect 146944 631518 146996 631524
rect 142816 631446 142844 631518
rect 146956 631446 146984 631518
rect 142804 631440 142856 631446
rect 101770 631408 101826 631417
rect 101476 631366 101770 631394
rect 143264 631440 143316 631446
rect 142804 631382 142856 631388
rect 142968 631388 143264 631394
rect 142968 631382 143316 631388
rect 146944 631440 146996 631446
rect 169668 631440 169720 631446
rect 146944 631382 146996 631388
rect 169372 631388 169668 631394
rect 188528 631440 188580 631446
rect 169372 631382 169720 631388
rect 188232 631388 188528 631394
rect 211068 631440 211120 631446
rect 188232 631382 188580 631388
rect 210864 631388 211068 631394
rect 233792 631440 233844 631446
rect 210864 631382 211120 631388
rect 233496 631388 233792 631394
rect 366560 631417 366588 634238
rect 369320 631938 369348 638250
rect 403256 638172 403308 638178
rect 403256 638114 403308 638120
rect 388168 637832 388220 637838
rect 388168 637774 388220 637780
rect 372712 635316 372764 635322
rect 372712 635258 372764 635264
rect 369288 631910 369348 631938
rect 372724 631938 372752 635258
rect 384028 635180 384080 635186
rect 384028 635122 384080 635128
rect 376852 632596 376904 632602
rect 376852 632538 376904 632544
rect 372724 631910 373060 631938
rect 376864 631802 376892 632538
rect 380256 632392 380308 632398
rect 380256 632334 380308 632340
rect 380268 631938 380296 632334
rect 384040 631938 384068 635122
rect 388180 631938 388208 637774
rect 395344 635044 395396 635050
rect 395344 634986 395396 634992
rect 391940 633888 391992 633894
rect 391940 633830 391992 633836
rect 391952 631938 391980 633830
rect 380268 631910 380604 631938
rect 384040 631910 384376 631938
rect 388148 631910 388208 631938
rect 391920 631910 391980 631938
rect 395356 631938 395384 634986
rect 399116 632256 399168 632262
rect 399116 632198 399168 632204
rect 399128 631938 399156 632198
rect 403268 631938 403296 638114
rect 422116 637968 422168 637974
rect 422116 637910 422168 637916
rect 410432 637764 410484 637770
rect 410432 637706 410484 637712
rect 406660 634976 406712 634982
rect 406660 634918 406712 634924
rect 395356 631910 395692 631938
rect 399128 631910 399464 631938
rect 403236 631910 403296 631938
rect 406672 631938 406700 634918
rect 410444 631938 410472 637706
rect 414204 636880 414256 636886
rect 414204 636822 414256 636828
rect 414216 631938 414244 636822
rect 422128 631938 422156 637910
rect 429212 635594 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 639606 462360 703520
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 462320 639600 462372 639606
rect 462320 639542 462372 639548
rect 440608 636744 440660 636750
rect 440608 636686 440660 636692
rect 429200 635588 429252 635594
rect 429200 635530 429252 635536
rect 433432 634364 433484 634370
rect 433432 634306 433484 634312
rect 425520 633820 425572 633826
rect 425520 633762 425572 633768
rect 406672 631910 407008 631938
rect 410444 631910 410780 631938
rect 414216 631910 414552 631938
rect 422096 631910 422156 631938
rect 425532 631938 425560 633762
rect 425532 631910 425868 631938
rect 433444 631802 433472 634306
rect 436836 633752 436888 633758
rect 436836 633694 436888 633700
rect 436848 631938 436876 633694
rect 440620 631938 440648 636686
rect 463240 636608 463292 636614
rect 463240 636550 463292 636556
rect 451924 636336 451976 636342
rect 451924 636278 451976 636284
rect 448520 633684 448572 633690
rect 448520 633626 448572 633632
rect 444702 632188 444754 632194
rect 444702 632130 444754 632136
rect 436848 631910 437184 631938
rect 440620 631910 440956 631938
rect 444714 631924 444742 632130
rect 448532 631938 448560 633626
rect 448500 631910 448560 631938
rect 451936 631938 451964 636278
rect 459560 634296 459612 634302
rect 459560 634238 459612 634244
rect 455696 633616 455748 633622
rect 455696 633558 455748 633564
rect 455708 631938 455736 633558
rect 459572 631938 459600 634238
rect 463252 631938 463280 636550
rect 474740 636540 474792 636546
rect 474740 636482 474792 636488
rect 470876 633548 470928 633554
rect 470876 633490 470928 633496
rect 467332 632224 467388 632233
rect 467332 632159 467388 632168
rect 451936 631910 452272 631938
rect 455708 631910 456044 631938
rect 459572 631910 459816 631938
rect 463252 631910 463588 631938
rect 467346 631924 467374 632159
rect 470888 631938 470916 633490
rect 474752 631938 474780 636482
rect 485872 636472 485924 636478
rect 485872 636414 485924 636420
rect 478326 633992 478382 634001
rect 478326 633927 478382 633936
rect 478340 631938 478368 633927
rect 482100 633480 482152 633486
rect 482100 633422 482152 633428
rect 482112 631938 482140 633422
rect 485884 631938 485912 636414
rect 494072 635526 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 638382 527220 703520
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700330 559696 703520
rect 549904 700324 549956 700330
rect 549904 700266 549956 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 527180 638376 527232 638382
rect 527180 638318 527232 638324
rect 522396 638240 522448 638246
rect 522396 638182 522448 638188
rect 521016 638104 521068 638110
rect 521016 638046 521068 638052
rect 520924 638036 520976 638042
rect 520924 637978 520976 637984
rect 518256 637900 518308 637906
rect 518256 637842 518308 637848
rect 515404 637696 515456 637702
rect 515404 637638 515456 637644
rect 514208 636676 514260 636682
rect 514208 636618 514260 636624
rect 497188 636404 497240 636410
rect 497188 636346 497240 636352
rect 494060 635520 494112 635526
rect 494060 635462 494112 635468
rect 490010 633720 490066 633729
rect 490010 633655 490066 633664
rect 470888 631910 471132 631938
rect 474752 631910 474904 631938
rect 478340 631910 478676 631938
rect 482112 631910 482448 631938
rect 485884 631910 486220 631938
rect 490024 631802 490052 633655
rect 493968 633480 494020 633486
rect 493968 633422 494020 633428
rect 493980 631938 494008 633422
rect 493764 631910 494008 631938
rect 497200 631938 497228 636346
rect 514022 636304 514078 636313
rect 514022 636239 514078 636248
rect 512828 635452 512880 635458
rect 512828 635394 512880 635400
rect 512736 635384 512788 635390
rect 512736 635326 512788 635332
rect 512642 634944 512698 634953
rect 512642 634879 512698 634888
rect 505376 633616 505428 633622
rect 505376 633558 505428 633564
rect 512000 633616 512052 633622
rect 512000 633558 512052 633564
rect 501604 633548 501656 633554
rect 501604 633490 501656 633496
rect 501616 631938 501644 633490
rect 505388 631938 505416 633558
rect 511080 633548 511132 633554
rect 511080 633490 511132 633496
rect 497200 631910 497536 631938
rect 501308 631910 501644 631938
rect 505080 631910 505416 631938
rect 376832 631774 376892 631802
rect 433412 631774 433472 631802
rect 489992 631774 490052 631802
rect 410064 631712 410116 631718
rect 410064 631654 410116 631660
rect 421012 631712 421064 631718
rect 421012 631654 421064 631660
rect 410076 631446 410104 631654
rect 415490 631544 415546 631553
rect 415490 631479 415546 631488
rect 416594 631544 416650 631553
rect 421024 631514 421052 631654
rect 416594 631479 416650 631488
rect 421012 631508 421064 631514
rect 415504 631446 415532 631479
rect 416608 631446 416636 631479
rect 421012 631450 421064 631456
rect 410064 631440 410116 631446
rect 233496 631382 233844 631388
rect 366546 631408 366602 631417
rect 142968 631366 143304 631382
rect 169372 631366 169708 631382
rect 188232 631366 188568 631382
rect 210864 631366 211108 631382
rect 233496 631366 233832 631382
rect 101770 631343 101826 631352
rect 410524 631440 410576 631446
rect 410064 631382 410116 631388
rect 410522 631408 410524 631417
rect 415492 631440 415544 631446
rect 410576 631408 410578 631417
rect 366546 631343 366602 631352
rect 415492 631382 415544 631388
rect 416596 631440 416648 631446
rect 429292 631440 429344 631446
rect 416596 631382 416648 631388
rect 417974 631408 418030 631417
rect 410522 631343 410578 631352
rect 418030 631366 418324 631394
rect 429344 631388 429640 631394
rect 429292 631382 429640 631388
rect 429304 631366 429640 631382
rect 417974 631343 418030 631352
rect 88306 71890 88334 72148
rect 89134 71890 89162 72148
rect 88306 71862 88380 71890
rect 77300 70236 77352 70242
rect 77300 70178 77352 70184
rect 74540 58744 74592 58750
rect 74540 58686 74592 58692
rect 72424 33108 72476 33114
rect 72424 33050 72476 33056
rect 73160 26920 73212 26926
rect 73160 26862 73212 26868
rect 73172 16574 73200 26862
rect 74552 16574 74580 58686
rect 77312 16574 77340 70178
rect 80060 66972 80112 66978
rect 80060 66914 80112 66920
rect 80072 16574 80100 66914
rect 88352 66910 88380 71862
rect 89088 71862 89162 71890
rect 89720 71936 89772 71942
rect 89962 71890 89990 72148
rect 90790 71942 90818 72148
rect 89720 71878 89772 71884
rect 89088 68338 89116 71862
rect 89076 68332 89128 68338
rect 89076 68274 89128 68280
rect 88340 66904 88392 66910
rect 88340 66846 88392 66852
rect 84200 64252 84252 64258
rect 84200 64194 84252 64200
rect 70412 16546 71544 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 77312 16546 78168 16574
rect 80072 16546 80928 16574
rect 69112 14476 69164 14482
rect 69112 14418 69164 14424
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 69124 480 69152 14418
rect 69940 3392 69992 3398
rect 69940 3334 69992 3340
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3334
rect 71516 480 71544 16546
rect 72608 5024 72660 5030
rect 72608 4966 72660 4972
rect 72620 480 72648 4966
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 77392 6656 77444 6662
rect 77392 6598 77444 6604
rect 76196 5092 76248 5098
rect 76196 5034 76248 5040
rect 76208 480 76236 5034
rect 77404 480 77432 6598
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 79692 5160 79744 5166
rect 79692 5102 79744 5108
rect 79704 480 79732 5102
rect 80900 480 80928 16546
rect 83280 5228 83332 5234
rect 83280 5170 83332 5176
rect 82084 3800 82136 3806
rect 82084 3742 82136 3748
rect 82096 480 82124 3742
rect 83292 480 83320 5170
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 64194
rect 85580 38004 85632 38010
rect 85580 37946 85632 37952
rect 85592 16574 85620 37946
rect 86960 28280 87012 28286
rect 86960 28222 87012 28228
rect 86972 16574 87000 28222
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 85684 480 85712 16546
rect 86868 5296 86920 5302
rect 86868 5238 86920 5244
rect 86880 480 86908 5238
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89732 6186 89760 71878
rect 89824 71862 89990 71890
rect 90778 71936 90830 71942
rect 91618 71890 91646 72148
rect 90778 71878 90830 71884
rect 91572 71862 91646 71890
rect 92446 71890 92474 72148
rect 93274 71890 93302 72148
rect 94102 71890 94130 72148
rect 94930 71890 94958 72148
rect 95758 71890 95786 72148
rect 92446 71862 92520 71890
rect 89824 42090 89852 71862
rect 91572 69698 91600 71862
rect 91560 69692 91612 69698
rect 91560 69634 91612 69640
rect 89812 42084 89864 42090
rect 89812 42026 89864 42032
rect 91100 31068 91152 31074
rect 91100 31010 91152 31016
rect 91112 16574 91140 31010
rect 91112 16546 91600 16574
rect 89720 6180 89772 6186
rect 89720 6122 89772 6128
rect 90364 5364 90416 5370
rect 90364 5306 90416 5312
rect 89168 3868 89220 3874
rect 89168 3810 89220 3816
rect 89180 480 89208 3810
rect 90376 480 90404 5306
rect 91572 480 91600 16546
rect 92492 3466 92520 71862
rect 92584 71862 93302 71890
rect 93964 71862 94130 71890
rect 94240 71862 94958 71890
rect 95712 71862 95786 71890
rect 96586 71890 96614 72148
rect 97414 71890 97442 72148
rect 98242 71890 98270 72148
rect 99070 71890 99098 72148
rect 99898 71890 99926 72148
rect 96586 71862 96660 71890
rect 92584 7614 92612 71862
rect 93860 68332 93912 68338
rect 93860 68274 93912 68280
rect 92664 49088 92716 49094
rect 92664 49030 92716 49036
rect 92676 16574 92704 49030
rect 92676 16546 92796 16574
rect 92572 7608 92624 7614
rect 92572 7550 92624 7556
rect 92480 3460 92532 3466
rect 92480 3402 92532 3408
rect 92768 480 92796 16546
rect 93872 5522 93900 68274
rect 93964 6254 93992 71862
rect 94240 60042 94268 71862
rect 95712 69766 95740 71862
rect 95700 69760 95752 69766
rect 95700 69702 95752 69708
rect 94228 60036 94280 60042
rect 94228 59978 94280 59984
rect 93952 6248 94004 6254
rect 93952 6190 94004 6196
rect 93872 5494 94728 5522
rect 93952 5432 94004 5438
rect 93952 5374 94004 5380
rect 93964 480 93992 5374
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 354 94728 5494
rect 96632 4826 96660 71862
rect 96724 71862 97442 71890
rect 98012 71862 98270 71890
rect 98656 71862 99098 71890
rect 99392 71862 99926 71890
rect 100726 71890 100754 72148
rect 101554 71890 101582 72148
rect 102382 71890 102410 72148
rect 103210 71890 103238 72148
rect 104038 71890 104066 72148
rect 100726 71862 100800 71890
rect 96724 43450 96752 71862
rect 96712 43444 96764 43450
rect 96712 43386 96764 43392
rect 96620 4820 96672 4826
rect 96620 4762 96672 4768
rect 97448 4820 97500 4826
rect 97448 4762 97500 4768
rect 96252 3460 96304 3466
rect 96252 3402 96304 3408
rect 96264 480 96292 3402
rect 97460 480 97488 4762
rect 98012 3534 98040 71862
rect 98656 64874 98684 71862
rect 98104 64846 98684 64874
rect 98104 3602 98132 64846
rect 98184 35216 98236 35222
rect 98184 35158 98236 35164
rect 98092 3596 98144 3602
rect 98092 3538 98144 3544
rect 98000 3528 98052 3534
rect 98000 3470 98052 3476
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 35158
rect 99392 4894 99420 71862
rect 100772 57254 100800 71862
rect 101508 71862 101582 71890
rect 102336 71862 102410 71890
rect 102520 71862 103238 71890
rect 103532 71862 104066 71890
rect 104866 71890 104894 72148
rect 105694 71890 105722 72148
rect 106522 71890 106550 72148
rect 107350 71890 107378 72148
rect 108178 71890 108206 72148
rect 104866 71862 104940 71890
rect 101508 69834 101536 71862
rect 102336 69970 102364 71862
rect 102324 69964 102376 69970
rect 102324 69906 102376 69912
rect 101496 69828 101548 69834
rect 101496 69770 101548 69776
rect 100760 57248 100812 57254
rect 100760 57190 100812 57196
rect 102232 50448 102284 50454
rect 102232 50390 102284 50396
rect 99472 40792 99524 40798
rect 99472 40734 99524 40740
rect 99484 16574 99512 40734
rect 100760 18624 100812 18630
rect 100760 18566 100812 18572
rect 99484 16546 99880 16574
rect 99380 4888 99432 4894
rect 99380 4830 99432 4836
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 18566
rect 102244 480 102272 50390
rect 102324 42084 102376 42090
rect 102324 42026 102376 42032
rect 102336 16574 102364 42026
rect 102336 16546 102456 16574
rect 102428 3482 102456 16546
rect 102520 4962 102548 71862
rect 103532 21418 103560 71862
rect 104912 69086 104940 71862
rect 105004 71862 105722 71890
rect 106384 71862 106550 71890
rect 106660 71862 107378 71890
rect 108132 71862 108206 71890
rect 109006 71890 109034 72148
rect 109834 71890 109862 72148
rect 109006 71862 109080 71890
rect 104164 69080 104216 69086
rect 104164 69022 104216 69028
rect 104900 69080 104952 69086
rect 104900 69022 104952 69028
rect 103520 21412 103572 21418
rect 103520 21354 103572 21360
rect 103612 21412 103664 21418
rect 103612 21354 103664 21360
rect 103624 16574 103652 21354
rect 103624 16546 104112 16574
rect 102508 4956 102560 4962
rect 102508 4898 102560 4904
rect 102428 3454 103376 3482
rect 103348 480 103376 3454
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 104176 11762 104204 69022
rect 105004 50386 105032 71862
rect 106280 69692 106332 69698
rect 106280 69634 106332 69640
rect 104992 50380 105044 50386
rect 104992 50322 105044 50328
rect 106292 16574 106320 69634
rect 106384 36582 106412 71862
rect 106660 58682 106688 71862
rect 108132 69902 108160 71862
rect 108120 69896 108172 69902
rect 108120 69838 108172 69844
rect 109052 64190 109080 71862
rect 109236 71862 109862 71890
rect 110420 71936 110472 71942
rect 110662 71890 110690 72148
rect 111490 71942 111518 72148
rect 110420 71878 110472 71884
rect 109040 64184 109092 64190
rect 109040 64126 109092 64132
rect 106648 58676 106700 58682
rect 106648 58618 106700 58624
rect 109236 55894 109264 71862
rect 109224 55888 109276 55894
rect 109224 55830 109276 55836
rect 106372 36576 106424 36582
rect 106372 36518 106424 36524
rect 107660 32428 107712 32434
rect 107660 32370 107712 32376
rect 107672 16574 107700 32370
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 104164 11756 104216 11762
rect 104164 11698 104216 11704
rect 105728 7608 105780 7614
rect 105728 7550 105780 7556
rect 105740 480 105768 7550
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 9036 109368 9042
rect 109316 8978 109368 8984
rect 109328 480 109356 8978
rect 110432 8974 110460 71878
rect 110616 71862 110690 71890
rect 111478 71936 111530 71942
rect 112318 71890 112346 72148
rect 111478 71878 111530 71884
rect 111904 71862 112346 71890
rect 113146 71890 113174 72148
rect 113974 71890 114002 72148
rect 113146 71862 113220 71890
rect 110512 44940 110564 44946
rect 110512 44882 110564 44888
rect 110420 8968 110472 8974
rect 110420 8910 110472 8916
rect 110524 480 110552 44882
rect 110616 33794 110644 71862
rect 111800 39500 111852 39506
rect 111800 39442 111852 39448
rect 110604 33788 110656 33794
rect 110604 33730 110656 33736
rect 111812 16574 111840 39442
rect 111904 39370 111932 71862
rect 113192 70038 113220 71862
rect 113284 71862 114002 71890
rect 114560 71936 114612 71942
rect 114802 71890 114830 72148
rect 115630 71942 115658 72148
rect 114560 71878 114612 71884
rect 113180 70032 113232 70038
rect 113180 69974 113232 69980
rect 111892 39364 111944 39370
rect 111892 39306 111944 39312
rect 113284 37942 113312 71862
rect 113272 37936 113324 37942
rect 113272 37878 113324 37884
rect 111812 16546 112392 16574
rect 111616 10396 111668 10402
rect 111616 10338 111668 10344
rect 111628 480 111656 10338
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 3936 114060 3942
rect 114008 3878 114060 3884
rect 114020 480 114048 3878
rect 114572 3670 114600 71878
rect 114664 71862 114830 71890
rect 115618 71936 115670 71942
rect 116458 71890 116486 72148
rect 115618 71878 115670 71884
rect 116044 71862 116486 71890
rect 117286 71890 117314 72148
rect 118114 71890 118142 72148
rect 118942 72026 118970 72148
rect 117286 71862 117360 71890
rect 114664 51746 114692 71862
rect 115940 66904 115992 66910
rect 115940 66846 115992 66852
rect 114652 51740 114704 51746
rect 114652 51682 114704 51688
rect 114652 33788 114704 33794
rect 114652 33730 114704 33736
rect 114664 16574 114692 33730
rect 115952 16574 115980 66846
rect 116044 22778 116072 71862
rect 117332 53106 117360 71862
rect 118068 71862 118142 71890
rect 118896 71998 118970 72026
rect 118068 70174 118096 71862
rect 118056 70168 118108 70174
rect 118056 70110 118108 70116
rect 117964 69080 118016 69086
rect 117964 69022 118016 69028
rect 117320 53100 117372 53106
rect 117320 53042 117372 53048
rect 116032 22772 116084 22778
rect 116032 22714 116084 22720
rect 114664 16546 114784 16574
rect 115952 16546 116440 16574
rect 114560 3664 114612 3670
rect 114560 3606 114612 3612
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117976 3738 118004 69022
rect 118896 65550 118924 71998
rect 119770 71890 119798 72148
rect 120598 71890 120626 72148
rect 119264 71862 119798 71890
rect 120552 71862 120626 71890
rect 121426 71890 121454 72148
rect 122254 71890 122282 72148
rect 121426 71862 121684 71890
rect 118884 65544 118936 65550
rect 118884 65486 118936 65492
rect 119264 64874 119292 71862
rect 120552 69086 120580 71862
rect 120540 69080 120592 69086
rect 120540 69022 120592 69028
rect 118712 64846 119292 64874
rect 118712 54534 118740 64846
rect 121552 62960 121604 62966
rect 121552 62902 121604 62908
rect 118700 54528 118752 54534
rect 118700 54470 118752 54476
rect 118700 36576 118752 36582
rect 118700 36518 118752 36524
rect 117964 3732 118016 3738
rect 117964 3674 118016 3680
rect 117596 3596 117648 3602
rect 117596 3538 117648 3544
rect 117608 480 117636 3538
rect 118712 3534 118740 36518
rect 121564 16574 121592 62902
rect 121656 62830 121684 71862
rect 121748 71862 122282 71890
rect 122840 71936 122892 71942
rect 123082 71890 123110 72148
rect 123910 71942 123938 72148
rect 122840 71878 122892 71884
rect 121644 62824 121696 62830
rect 121644 62766 121696 62772
rect 121564 16546 121684 16574
rect 118792 6180 118844 6186
rect 118792 6122 118844 6128
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 118804 480 118832 6122
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 121092 3528 121144 3534
rect 121092 3470 121144 3476
rect 121656 3482 121684 16546
rect 121748 6322 121776 71862
rect 122852 15910 122880 71878
rect 122944 71862 123110 71890
rect 123898 71936 123950 71942
rect 124738 71890 124766 72148
rect 123898 71878 123950 71884
rect 124324 71862 124766 71890
rect 125566 71890 125594 72148
rect 126394 71890 126422 72148
rect 127222 71890 127250 72148
rect 128050 71890 128078 72148
rect 128878 71890 128906 72148
rect 125566 71862 125640 71890
rect 122944 49026 122972 71862
rect 124220 69760 124272 69766
rect 124220 69702 124272 69708
rect 122932 49020 122984 49026
rect 122932 48962 122984 48968
rect 122840 15904 122892 15910
rect 122840 15846 122892 15852
rect 123024 15904 123076 15910
rect 123024 15846 123076 15852
rect 121736 6316 121788 6322
rect 121736 6258 121788 6264
rect 119908 480 119936 3470
rect 121104 480 121132 3470
rect 121656 3454 122328 3482
rect 122300 480 122328 3454
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 15846
rect 124232 1306 124260 69702
rect 124324 6390 124352 71862
rect 125612 40730 125640 71862
rect 125704 71862 126422 71890
rect 126992 71862 127250 71890
rect 127544 71862 128078 71890
rect 128372 71862 128906 71890
rect 129706 71890 129734 72148
rect 130534 71890 130562 72148
rect 129706 71862 129780 71890
rect 125704 44878 125732 71862
rect 125692 44872 125744 44878
rect 125692 44814 125744 44820
rect 125600 40724 125652 40730
rect 125600 40666 125652 40672
rect 126992 24138 127020 71862
rect 127544 64874 127572 71862
rect 127084 64846 127572 64874
rect 127084 42158 127112 64846
rect 127072 42152 127124 42158
rect 127072 42094 127124 42100
rect 126980 24132 127032 24138
rect 126980 24074 127032 24080
rect 127072 24132 127124 24138
rect 127072 24074 127124 24080
rect 125876 7676 125928 7682
rect 125876 7618 125928 7624
rect 124312 6384 124364 6390
rect 124312 6326 124364 6332
rect 124232 1278 124720 1306
rect 124692 480 124720 1278
rect 125888 480 125916 7618
rect 127084 6914 127112 24074
rect 128372 17270 128400 71862
rect 128360 17264 128412 17270
rect 128360 17206 128412 17212
rect 128912 11756 128964 11762
rect 128912 11698 128964 11704
rect 128176 8968 128228 8974
rect 128176 8910 128228 8916
rect 126992 6886 127112 6914
rect 126992 480 127020 6886
rect 128188 480 128216 8910
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 11698
rect 129752 6458 129780 71862
rect 129844 71862 130562 71890
rect 131120 71936 131172 71942
rect 131362 71890 131390 72148
rect 132190 71942 132218 72148
rect 131120 71878 131172 71884
rect 129844 29646 129872 71862
rect 129832 29640 129884 29646
rect 129832 29582 129884 29588
rect 129832 22772 129884 22778
rect 129832 22714 129884 22720
rect 129844 16574 129872 22714
rect 129844 16546 130608 16574
rect 129740 6452 129792 6458
rect 129740 6394 129792 6400
rect 130580 480 130608 16546
rect 131132 6526 131160 71878
rect 131224 71862 131390 71890
rect 132178 71936 132230 71942
rect 133018 71890 133046 72148
rect 132178 71878 132230 71884
rect 132512 71862 133046 71890
rect 133846 71890 133874 72148
rect 134674 71890 134702 72148
rect 133846 71862 133920 71890
rect 131224 46238 131252 71862
rect 131212 46232 131264 46238
rect 131212 46174 131264 46180
rect 132512 43518 132540 71862
rect 132500 43512 132552 43518
rect 132500 43454 132552 43460
rect 132960 13116 133012 13122
rect 132960 13058 133012 13064
rect 131120 6520 131172 6526
rect 131120 6462 131172 6468
rect 131764 6248 131816 6254
rect 131764 6190 131816 6196
rect 131776 480 131804 6190
rect 132972 480 133000 13058
rect 133892 10334 133920 71862
rect 134168 71862 134702 71890
rect 135260 71936 135312 71942
rect 135502 71890 135530 72148
rect 136330 71942 136358 72148
rect 135260 71878 135312 71884
rect 134064 25628 134116 25634
rect 134064 25570 134116 25576
rect 133880 10328 133932 10334
rect 133880 10270 133932 10276
rect 134076 1442 134104 25570
rect 134168 6594 134196 71862
rect 135272 14482 135300 71878
rect 135364 71862 135530 71890
rect 136318 71936 136370 71942
rect 137158 71890 137186 72148
rect 136318 71878 136370 71884
rect 136652 71862 137186 71890
rect 137986 71890 138014 72148
rect 138814 71890 138842 72148
rect 139642 71890 139670 72148
rect 140470 71890 140498 72148
rect 141298 71890 141326 72148
rect 137986 71862 138060 71890
rect 135364 57322 135392 71862
rect 135904 69964 135956 69970
rect 135904 69906 135956 69912
rect 135352 57316 135404 57322
rect 135352 57258 135404 57264
rect 135352 29640 135404 29646
rect 135352 29582 135404 29588
rect 135260 14476 135312 14482
rect 135260 14418 135312 14424
rect 135364 6914 135392 29582
rect 135812 14476 135864 14482
rect 135812 14418 135864 14424
rect 135272 6886 135392 6914
rect 134156 6588 134208 6594
rect 134156 6530 134208 6536
rect 134076 1414 134196 1442
rect 134168 480 134196 1414
rect 135272 480 135300 6886
rect 135824 3482 135852 14418
rect 135916 3806 135944 69906
rect 136652 25566 136680 71862
rect 138032 70106 138060 71862
rect 138216 71862 138842 71890
rect 139412 71862 139670 71890
rect 139872 71862 140498 71890
rect 140792 71862 141326 71890
rect 142126 71890 142154 72148
rect 142954 71890 142982 72148
rect 143782 71890 143810 72148
rect 144610 71890 144638 72148
rect 145438 71890 145466 72148
rect 142126 71862 142200 71890
rect 138020 70100 138072 70106
rect 138020 70042 138072 70048
rect 136640 25560 136692 25566
rect 136640 25502 136692 25508
rect 137192 11824 137244 11830
rect 137192 11766 137244 11772
rect 135904 3800 135956 3806
rect 135904 3742 135956 3748
rect 135824 3454 136496 3482
rect 136468 480 136496 3454
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 11766
rect 138216 5030 138244 71862
rect 139412 26926 139440 71862
rect 139872 64874 139900 71862
rect 140044 69896 140096 69902
rect 140044 69838 140096 69844
rect 139504 64846 139900 64874
rect 139504 58750 139532 64846
rect 139492 58744 139544 58750
rect 139492 58686 139544 58692
rect 139400 26920 139452 26926
rect 139400 26862 139452 26868
rect 139584 15972 139636 15978
rect 139584 15914 139636 15920
rect 138848 6316 138900 6322
rect 138848 6258 138900 6264
rect 138204 5024 138256 5030
rect 138204 4966 138256 4972
rect 138860 480 138888 6258
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 15914
rect 140056 3874 140084 69838
rect 140792 5098 140820 71862
rect 142172 6662 142200 71862
rect 142908 71862 142982 71890
rect 143552 71862 143810 71890
rect 144564 71862 144638 71890
rect 145392 71862 145466 71890
rect 146266 71890 146294 72148
rect 147094 71890 147122 72148
rect 146266 71862 146340 71890
rect 142908 70242 142936 71862
rect 142896 70236 142948 70242
rect 142896 70178 142948 70184
rect 142252 43444 142304 43450
rect 142252 43386 142304 43392
rect 142160 6656 142212 6662
rect 142160 6598 142212 6604
rect 140780 5092 140832 5098
rect 140780 5034 140832 5040
rect 141240 4888 141292 4894
rect 141240 4830 141292 4836
rect 140044 3868 140096 3874
rect 140044 3810 140096 3816
rect 141252 480 141280 4830
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142264 354 142292 43386
rect 143552 6914 143580 71862
rect 144184 69828 144236 69834
rect 144184 69770 144236 69776
rect 143632 17264 143684 17270
rect 143632 17206 143684 17212
rect 143644 16574 143672 17206
rect 143644 16546 143764 16574
rect 143552 6886 143672 6914
rect 143644 5166 143672 6886
rect 143632 5160 143684 5166
rect 143632 5102 143684 5108
rect 143736 3482 143764 16546
rect 143552 3454 143764 3482
rect 144196 3466 144224 69770
rect 144564 66978 144592 71862
rect 145392 69970 145420 71862
rect 145380 69964 145432 69970
rect 145380 69906 145432 69912
rect 144552 66972 144604 66978
rect 144552 66914 144604 66920
rect 144920 55888 144972 55894
rect 144920 55830 144972 55836
rect 144932 16574 144960 55830
rect 144932 16546 145512 16574
rect 144736 4956 144788 4962
rect 144736 4898 144788 4904
rect 144184 3460 144236 3466
rect 143552 480 143580 3454
rect 144184 3402 144236 3408
rect 144748 480 144776 4898
rect 142406 354 142518 480
rect 142264 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146312 5234 146340 71862
rect 146496 71862 147122 71890
rect 147680 71936 147732 71942
rect 147922 71890 147950 72148
rect 148750 71942 148778 72148
rect 147680 71878 147732 71884
rect 146392 64388 146444 64394
rect 146392 64330 146444 64336
rect 146404 16574 146432 64330
rect 146496 64258 146524 71862
rect 146484 64252 146536 64258
rect 146484 64194 146536 64200
rect 146404 16546 147168 16574
rect 146300 5228 146352 5234
rect 146300 5170 146352 5176
rect 147140 480 147168 16546
rect 147692 5302 147720 71878
rect 147784 71862 147950 71890
rect 148738 71936 148790 71942
rect 149578 71890 149606 72148
rect 148738 71878 148790 71884
rect 149164 71862 149606 71890
rect 150406 71890 150434 72148
rect 151234 71890 151262 72148
rect 152062 71890 152090 72148
rect 152890 71890 152918 72148
rect 153718 71890 153746 72148
rect 150406 71862 150480 71890
rect 147784 38010 147812 71862
rect 149060 68400 149112 68406
rect 149060 68342 149112 68348
rect 147772 38004 147824 38010
rect 147772 37946 147824 37952
rect 147772 26920 147824 26926
rect 147772 26862 147824 26868
rect 147784 16574 147812 26862
rect 149072 16574 149100 68342
rect 149164 28286 149192 71862
rect 150452 69902 150480 71862
rect 150636 71862 151262 71890
rect 151924 71862 152090 71890
rect 152200 71862 152918 71890
rect 153212 71862 153746 71890
rect 154546 71890 154574 72148
rect 155374 71890 155402 72148
rect 156202 71890 156230 72148
rect 157030 71890 157058 72148
rect 157858 71890 157886 72148
rect 154546 71862 154620 71890
rect 150440 69896 150492 69902
rect 150440 69838 150492 69844
rect 149152 28280 149204 28286
rect 149152 28222 149204 28228
rect 150636 16574 150664 71862
rect 151820 51740 151872 51746
rect 151820 51682 151872 51688
rect 147784 16546 147904 16574
rect 149072 16546 149560 16574
rect 150636 16546 150756 16574
rect 147680 5296 147732 5302
rect 147680 5238 147732 5244
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150624 13184 150676 13190
rect 150624 13126 150676 13132
rect 150636 480 150664 13126
rect 150728 5370 150756 16546
rect 151832 9674 151860 51682
rect 151924 31074 151952 71862
rect 152200 49094 152228 71862
rect 152188 49088 152240 49094
rect 152188 49030 152240 49036
rect 151912 31068 151964 31074
rect 151912 31010 151964 31016
rect 151912 28280 151964 28286
rect 151912 28222 151964 28228
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 28222
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 150716 5364 150768 5370
rect 150716 5306 150768 5312
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 153212 5438 153240 71862
rect 154592 68338 154620 71862
rect 155328 71862 155402 71890
rect 155972 71862 156230 71890
rect 156432 71862 157058 71890
rect 157352 71862 157886 71890
rect 158686 71890 158714 72148
rect 159514 71890 159542 72148
rect 158686 71862 158760 71890
rect 155328 69834 155356 71862
rect 155316 69828 155368 69834
rect 155316 69770 155368 69776
rect 154580 68332 154632 68338
rect 154580 68274 154632 68280
rect 153200 5432 153252 5438
rect 153200 5374 153252 5380
rect 154212 5024 154264 5030
rect 154212 4966 154264 4972
rect 154224 480 154252 4966
rect 155972 4826 156000 71862
rect 156432 64874 156460 71862
rect 156604 69828 156656 69834
rect 156604 69770 156656 69776
rect 156064 64846 156460 64874
rect 156064 35222 156092 64846
rect 156052 35216 156104 35222
rect 156052 35158 156104 35164
rect 156052 31068 156104 31074
rect 156052 31010 156104 31016
rect 156064 16574 156092 31010
rect 156064 16546 156184 16574
rect 155960 4820 156012 4826
rect 155960 4762 156012 4768
rect 155408 3052 155460 3058
rect 155408 2994 155460 3000
rect 155420 480 155448 2994
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 156616 3942 156644 69770
rect 157352 40798 157380 71862
rect 157984 65544 158036 65550
rect 157984 65486 158036 65492
rect 157340 40792 157392 40798
rect 157340 40734 157392 40740
rect 157340 18692 157392 18698
rect 157340 18634 157392 18640
rect 157352 16574 157380 18634
rect 157352 16546 157840 16574
rect 156604 3936 156656 3942
rect 156604 3878 156656 3884
rect 157812 480 157840 16546
rect 157996 3058 158024 65486
rect 158732 18630 158760 71862
rect 158824 71862 159542 71890
rect 160100 71936 160152 71942
rect 160342 71890 160370 72148
rect 161170 71942 161198 72148
rect 160100 71878 160152 71884
rect 158824 50454 158852 71862
rect 158812 50448 158864 50454
rect 158812 50390 158864 50396
rect 160112 21418 160140 71878
rect 160204 71862 160370 71890
rect 161158 71936 161210 71942
rect 161998 71890 162026 72148
rect 161158 71878 161210 71884
rect 161492 71862 162026 71890
rect 162826 71890 162854 72148
rect 163654 71890 163682 72148
rect 164482 71890 164510 72148
rect 165310 71890 165338 72148
rect 166138 71890 166166 72148
rect 162826 71862 162900 71890
rect 160204 42090 160232 71862
rect 160192 42084 160244 42090
rect 160192 42026 160244 42032
rect 160100 21412 160152 21418
rect 160100 21354 160152 21360
rect 158720 18624 158772 18630
rect 158720 18566 158772 18572
rect 158904 16040 158956 16046
rect 158904 15982 158956 15988
rect 157984 3052 158036 3058
rect 157984 2994 158036 3000
rect 158916 480 158944 15982
rect 161296 9104 161348 9110
rect 161296 9046 161348 9052
rect 160100 3460 160152 3466
rect 160100 3402 160152 3408
rect 160112 480 160140 3402
rect 161308 480 161336 9046
rect 161492 7614 161520 71862
rect 162872 69698 162900 71862
rect 162964 71862 163682 71890
rect 164436 71862 164510 71890
rect 165264 71862 165338 71890
rect 165724 71862 166166 71890
rect 166966 71890 166994 72148
rect 167794 71890 167822 72148
rect 168622 71890 168650 72148
rect 169450 71890 169478 72148
rect 170278 71890 170306 72148
rect 166966 71862 167040 71890
rect 162860 69692 162912 69698
rect 162860 69634 162912 69640
rect 162124 69080 162176 69086
rect 162124 69022 162176 69028
rect 162136 44946 162164 69022
rect 162124 44940 162176 44946
rect 162124 44882 162176 44888
rect 162964 32434 162992 71862
rect 162952 32428 163004 32434
rect 162952 32370 163004 32376
rect 161572 21412 161624 21418
rect 161572 21354 161624 21360
rect 161584 16574 161612 21354
rect 162860 17332 162912 17338
rect 162860 17274 162912 17280
rect 162872 16574 162900 17274
rect 164436 16574 164464 71862
rect 164884 69148 164936 69154
rect 164884 69090 164936 69096
rect 161584 16546 162072 16574
rect 162872 16546 163728 16574
rect 161480 7608 161532 7614
rect 161480 7550 161532 7556
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 164344 16546 164464 16574
rect 164344 9042 164372 16546
rect 164424 10328 164476 10334
rect 164424 10270 164476 10276
rect 164332 9036 164384 9042
rect 164332 8978 164384 8984
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 10270
rect 164896 3602 164924 69090
rect 165264 69086 165292 71862
rect 165252 69080 165304 69086
rect 165252 69022 165304 69028
rect 165620 66972 165672 66978
rect 165620 66914 165672 66920
rect 165632 6914 165660 66914
rect 165724 10402 165752 71862
rect 167012 39506 167040 71862
rect 167748 71862 167822 71890
rect 168392 71862 168650 71890
rect 169404 71862 169478 71890
rect 170232 71862 170306 71890
rect 171106 71890 171134 72148
rect 171934 71890 171962 72148
rect 172762 72026 172790 72148
rect 171106 71862 171272 71890
rect 167644 69896 167696 69902
rect 167644 69838 167696 69844
rect 167000 39500 167052 39506
rect 167000 39442 167052 39448
rect 165712 10396 165764 10402
rect 165712 10338 165764 10344
rect 165632 6886 166120 6914
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 166092 480 166120 6886
rect 167656 3534 167684 69838
rect 167748 69834 167776 71862
rect 167736 69828 167788 69834
rect 167736 69770 167788 69776
rect 168392 33794 168420 71862
rect 169404 66910 169432 71862
rect 169760 69692 169812 69698
rect 169760 69634 169812 69640
rect 169392 66904 169444 66910
rect 169392 66846 169444 66852
rect 168380 33788 168432 33794
rect 168380 33730 168432 33736
rect 169772 16574 169800 69634
rect 170232 69154 170260 71862
rect 170404 69828 170456 69834
rect 170404 69770 170456 69776
rect 170220 69148 170272 69154
rect 170220 69090 170272 69096
rect 169772 16546 170352 16574
rect 169576 9036 169628 9042
rect 169576 8978 169628 8984
rect 168380 7608 168432 7614
rect 168380 7550 168432 7556
rect 167644 3528 167696 3534
rect 167644 3470 167696 3476
rect 167184 3188 167236 3194
rect 167184 3130 167236 3136
rect 167196 480 167224 3130
rect 168392 480 168420 7550
rect 169588 480 169616 8978
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 170416 3194 170444 69770
rect 171140 68332 171192 68338
rect 171140 68274 171192 68280
rect 171152 3482 171180 68274
rect 171244 6186 171272 71862
rect 171336 71862 171962 71890
rect 172532 71998 172790 72026
rect 171336 36582 171364 71862
rect 172532 69902 172560 71998
rect 173590 71890 173618 72148
rect 174418 71890 174446 72148
rect 172624 71862 173618 71890
rect 173912 71862 174446 71890
rect 175246 71890 175274 72148
rect 176074 71890 176102 72148
rect 175246 71862 175320 71890
rect 172520 69896 172572 69902
rect 172520 69838 172572 69844
rect 172624 62966 172652 71862
rect 172612 62960 172664 62966
rect 172612 62902 172664 62908
rect 171324 36576 171376 36582
rect 171324 36518 171376 36524
rect 173912 15910 173940 71862
rect 174544 70032 174596 70038
rect 174544 69974 174596 69980
rect 173900 15904 173952 15910
rect 173900 15846 173952 15852
rect 171232 6180 171284 6186
rect 171232 6122 171284 6128
rect 173164 3528 173216 3534
rect 171152 3454 172008 3482
rect 173164 3470 173216 3476
rect 170404 3188 170456 3194
rect 170404 3130 170456 3136
rect 171980 480 172008 3454
rect 173176 480 173204 3470
rect 174268 3460 174320 3466
rect 174268 3402 174320 3408
rect 174280 480 174308 3402
rect 174556 3398 174584 69974
rect 175292 69766 175320 71862
rect 175384 71862 176102 71890
rect 176660 71936 176712 71942
rect 176902 71890 176930 72148
rect 177730 71942 177758 72148
rect 176660 71878 176712 71884
rect 175280 69760 175332 69766
rect 175280 69702 175332 69708
rect 175280 66904 175332 66910
rect 175280 66846 175332 66852
rect 174636 58676 174688 58682
rect 174636 58618 174688 58624
rect 174648 3534 174676 58618
rect 175292 6914 175320 66846
rect 175384 7682 175412 71862
rect 175924 21480 175976 21486
rect 175924 21422 175976 21428
rect 175372 7676 175424 7682
rect 175372 7618 175424 7624
rect 175292 6886 175504 6914
rect 174636 3528 174688 3534
rect 174636 3470 174688 3476
rect 174544 3392 174596 3398
rect 174544 3334 174596 3340
rect 175476 480 175504 6886
rect 175936 3466 175964 21422
rect 176672 8974 176700 71878
rect 176764 71862 176930 71890
rect 177718 71936 177770 71942
rect 178558 71890 178586 72148
rect 177718 71878 177770 71884
rect 178144 71862 178586 71890
rect 179386 71890 179414 72148
rect 180214 71890 180242 72148
rect 181042 71890 181070 72148
rect 181870 71890 181898 72148
rect 182698 71890 182726 72148
rect 179386 71862 179460 71890
rect 176764 24138 176792 71862
rect 178040 62824 178092 62830
rect 178040 62766 178092 62772
rect 176752 24132 176804 24138
rect 176752 24074 176804 24080
rect 176660 8968 176712 8974
rect 176660 8910 176712 8916
rect 178052 6914 178080 62766
rect 178144 11762 178172 71862
rect 179432 22778 179460 71862
rect 179616 71862 180242 71890
rect 180812 71862 181070 71890
rect 181456 71862 181898 71890
rect 182192 71862 182726 71890
rect 183526 71890 183554 72148
rect 184354 71890 184382 72148
rect 185182 71890 185210 72148
rect 186010 71890 186038 72148
rect 186838 71890 186866 72148
rect 183526 71862 183600 71890
rect 179420 22772 179472 22778
rect 179420 22714 179472 22720
rect 178132 11756 178184 11762
rect 178132 11698 178184 11704
rect 178684 10396 178736 10402
rect 178684 10338 178736 10344
rect 178052 6886 178632 6914
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 175924 3460 175976 3466
rect 175924 3402 175976 3408
rect 176672 480 176700 3470
rect 177856 3460 177908 3466
rect 177856 3402 177908 3408
rect 177868 480 177896 3402
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 6886
rect 178696 3534 178724 10338
rect 179616 6254 179644 71862
rect 180812 13122 180840 71862
rect 181456 64874 181484 71862
rect 180904 64846 181484 64874
rect 180904 25634 180932 64846
rect 182192 29646 182220 71862
rect 182824 57248 182876 57254
rect 182824 57190 182876 57196
rect 182180 29640 182232 29646
rect 182180 29582 182232 29588
rect 180892 25628 180944 25634
rect 180892 25570 180944 25576
rect 180800 13116 180852 13122
rect 180800 13058 180852 13064
rect 179604 6248 179656 6254
rect 179604 6190 179656 6196
rect 182548 6180 182600 6186
rect 182548 6122 182600 6128
rect 180248 4140 180300 4146
rect 180248 4082 180300 4088
rect 178684 3528 178736 3534
rect 178684 3470 178736 3476
rect 180260 480 180288 4082
rect 181444 3596 181496 3602
rect 181444 3538 181496 3544
rect 181456 480 181484 3538
rect 182560 480 182588 6122
rect 182836 4146 182864 57190
rect 183572 14482 183600 71862
rect 183848 71862 184382 71890
rect 185044 71862 185210 71890
rect 185320 71862 186038 71890
rect 186332 71862 186866 71890
rect 187666 71890 187694 72148
rect 188494 71890 188522 72148
rect 189322 71890 189350 72148
rect 190150 71890 190178 72148
rect 190978 71890 191006 72148
rect 187666 71862 187740 71890
rect 183560 14476 183612 14482
rect 183560 14418 183612 14424
rect 183744 14476 183796 14482
rect 183744 14418 183796 14424
rect 182824 4140 182876 4146
rect 182824 4082 182876 4088
rect 183756 480 183784 14418
rect 183848 11830 183876 71862
rect 184940 69760 184992 69766
rect 184940 69702 184992 69708
rect 183836 11824 183888 11830
rect 183836 11766 183888 11772
rect 184952 480 184980 69702
rect 185044 6322 185072 71862
rect 185320 15978 185348 71862
rect 185308 15972 185360 15978
rect 185308 15914 185360 15920
rect 186136 11756 186188 11762
rect 186136 11698 186188 11704
rect 185032 6316 185084 6322
rect 185032 6258 185084 6264
rect 186148 480 186176 11698
rect 186332 4894 186360 71862
rect 187712 43450 187740 71862
rect 187896 71862 188522 71890
rect 189092 71862 189350 71890
rect 189460 71862 190178 71890
rect 190472 71862 191006 71890
rect 191806 71890 191834 72148
rect 192634 71890 192662 72148
rect 193462 71890 193490 72148
rect 194290 71890 194318 72148
rect 195118 71890 195146 72148
rect 191806 71862 191972 71890
rect 187700 43444 187752 43450
rect 187700 43386 187752 43392
rect 187896 17270 187924 71862
rect 188344 50380 188396 50386
rect 188344 50322 188396 50328
rect 187884 17264 187936 17270
rect 187884 17206 187936 17212
rect 186320 4888 186372 4894
rect 186320 4830 186372 4836
rect 188356 3534 188384 50322
rect 189092 4962 189120 71862
rect 189172 64184 189224 64190
rect 189172 64126 189224 64132
rect 189184 16574 189212 64126
rect 189460 55894 189488 71862
rect 190472 64394 190500 71862
rect 191840 69896 191892 69902
rect 191840 69838 191892 69844
rect 190460 64388 190512 64394
rect 190460 64330 190512 64336
rect 189448 55888 189500 55894
rect 189448 55830 189500 55836
rect 191852 16574 191880 69838
rect 191944 26926 191972 71862
rect 192588 71862 192662 71890
rect 193324 71862 193490 71890
rect 193600 71862 194318 71890
rect 194612 71862 195146 71890
rect 195946 71890 195974 72148
rect 196774 71890 196802 72148
rect 195946 71862 196020 71890
rect 192588 68406 192616 71862
rect 192576 68400 192628 68406
rect 192576 68342 192628 68348
rect 193220 68400 193272 68406
rect 193220 68342 193272 68348
rect 192484 64252 192536 64258
rect 192484 64194 192536 64200
rect 191932 26920 191984 26926
rect 191932 26862 191984 26868
rect 189184 16546 189304 16574
rect 191852 16546 192064 16574
rect 189080 4956 189132 4962
rect 189080 4898 189132 4904
rect 188528 3596 188580 3602
rect 188528 3538 188580 3544
rect 187332 3528 187384 3534
rect 187332 3470 187384 3476
rect 188344 3528 188396 3534
rect 188344 3470 188396 3476
rect 187344 480 187372 3470
rect 188540 480 188568 3538
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 190840 480 190868 3334
rect 192036 480 192064 16546
rect 192496 3398 192524 64194
rect 192484 3392 192536 3398
rect 192484 3334 192536 3340
rect 193232 480 193260 68342
rect 193324 13190 193352 71862
rect 193600 28286 193628 71862
rect 194612 51746 194640 71862
rect 194600 51740 194652 51746
rect 194600 51682 194652 51688
rect 193588 28280 193640 28286
rect 193588 28222 193640 28228
rect 193312 13184 193364 13190
rect 193312 13126 193364 13132
rect 195992 5030 196020 71862
rect 196728 71862 196802 71890
rect 197452 71936 197504 71942
rect 197602 71890 197630 72148
rect 198430 71942 198458 72148
rect 197452 71878 197504 71884
rect 196072 65680 196124 65686
rect 196072 65622 196124 65628
rect 196084 16574 196112 65622
rect 196728 65550 196756 71862
rect 197360 69964 197412 69970
rect 197360 69906 197412 69912
rect 196716 65544 196768 65550
rect 196716 65486 196768 65492
rect 197372 16574 197400 69906
rect 197464 18698 197492 71878
rect 197556 71862 197630 71890
rect 198418 71936 198470 71942
rect 199258 71890 199286 72148
rect 198418 71878 198470 71884
rect 198844 71862 199286 71890
rect 200086 71890 200114 72148
rect 200914 71890 200942 72148
rect 200086 71862 200160 71890
rect 197556 31074 197584 71862
rect 198740 70100 198792 70106
rect 198740 70042 198792 70048
rect 197544 31068 197596 31074
rect 197544 31010 197596 31016
rect 197452 18692 197504 18698
rect 197452 18634 197504 18640
rect 196084 16546 196848 16574
rect 197372 16546 197952 16574
rect 195980 5024 196032 5030
rect 195980 4966 196032 4972
rect 194416 4820 194468 4826
rect 194416 4762 194468 4768
rect 194428 480 194456 4762
rect 195612 3664 195664 3670
rect 195612 3606 195664 3612
rect 195624 480 195652 3606
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 189694 -960 189806 326
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 70042
rect 198844 16046 198872 71862
rect 200132 70038 200160 71862
rect 200224 71862 200942 71890
rect 201500 71936 201552 71942
rect 201742 71890 201770 72148
rect 202570 71942 202598 72148
rect 201500 71878 201552 71884
rect 200120 70032 200172 70038
rect 200120 69974 200172 69980
rect 200120 67040 200172 67046
rect 200120 66982 200172 66988
rect 198832 16040 198884 16046
rect 198832 15982 198884 15988
rect 200132 6914 200160 66982
rect 200224 9110 200252 71862
rect 201512 17338 201540 71878
rect 201604 71862 201770 71890
rect 202558 71936 202610 71942
rect 203398 71890 203426 72148
rect 202558 71878 202610 71884
rect 202892 71862 203426 71890
rect 204226 71890 204254 72148
rect 205054 71890 205082 72148
rect 205882 71890 205910 72148
rect 206710 71890 206738 72148
rect 207538 71890 207566 72148
rect 204226 71862 204300 71890
rect 201604 21418 201632 71862
rect 201592 21412 201644 21418
rect 201592 21354 201644 21360
rect 201500 17332 201552 17338
rect 201500 17274 201552 17280
rect 202892 10334 202920 71862
rect 204272 66978 204300 71862
rect 205008 71862 205082 71890
rect 205744 71862 205910 71890
rect 206020 71862 206738 71890
rect 207492 71862 207566 71890
rect 208366 71890 208394 72148
rect 209194 71890 209222 72148
rect 210022 71890 210050 72148
rect 210850 71890 210878 72148
rect 211678 71890 211706 72148
rect 208366 71862 208440 71890
rect 205008 69834 205036 71862
rect 204996 69828 205048 69834
rect 204996 69770 205048 69776
rect 205640 69828 205692 69834
rect 205640 69770 205692 69776
rect 204260 66972 204312 66978
rect 204260 66914 204312 66920
rect 205088 13116 205140 13122
rect 205088 13058 205140 13064
rect 202880 10328 202932 10334
rect 202880 10270 202932 10276
rect 200212 9104 200264 9110
rect 200212 9046 200264 9052
rect 203892 7676 203944 7682
rect 203892 7618 203944 7624
rect 200132 6886 200344 6914
rect 200316 480 200344 6886
rect 201500 4004 201552 4010
rect 201500 3946 201552 3952
rect 201512 480 201540 3946
rect 202696 3732 202748 3738
rect 202696 3674 202748 3680
rect 202708 480 202736 3674
rect 203904 480 203932 7618
rect 205100 480 205128 13058
rect 205652 6914 205680 69770
rect 205744 7614 205772 71862
rect 206020 9042 206048 71862
rect 207492 69698 207520 71862
rect 207480 69692 207532 69698
rect 207480 69634 207532 69640
rect 207020 68468 207072 68474
rect 207020 68410 207072 68416
rect 206008 9036 206060 9042
rect 206008 8978 206060 8984
rect 205732 7608 205784 7614
rect 205732 7550 205784 7556
rect 205652 6886 206232 6914
rect 206204 480 206232 6886
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 68410
rect 208412 68338 208440 71862
rect 208596 71862 209222 71890
rect 209884 71862 210050 71890
rect 210804 71862 210878 71890
rect 211264 71862 211706 71890
rect 212506 71890 212534 72148
rect 213334 71890 213362 72148
rect 212506 71862 212580 71890
rect 208400 68332 208452 68338
rect 208400 68274 208452 68280
rect 208596 58682 208624 71862
rect 209780 67108 209832 67114
rect 209780 67050 209832 67056
rect 208584 58676 208636 58682
rect 208584 58618 208636 58624
rect 208584 4072 208636 4078
rect 208584 4014 208636 4020
rect 208596 480 208624 4014
rect 209792 3398 209820 67050
rect 209884 21486 209912 71862
rect 210424 69080 210476 69086
rect 210424 69022 210476 69028
rect 209872 21480 209924 21486
rect 209872 21422 209924 21428
rect 209872 3800 209924 3806
rect 209872 3742 209924 3748
rect 209780 3392 209832 3398
rect 209780 3334 209832 3340
rect 209884 1986 209912 3742
rect 210436 3466 210464 69022
rect 210804 66910 210832 71862
rect 210792 66904 210844 66910
rect 210792 66846 210844 66852
rect 211160 65544 211212 65550
rect 211160 65486 211212 65492
rect 211172 6914 211200 65486
rect 211264 10402 211292 71862
rect 212552 69086 212580 71862
rect 212644 71862 213362 71890
rect 213920 71936 213972 71942
rect 214162 71890 214190 72148
rect 214990 71942 215018 72148
rect 213920 71878 213972 71884
rect 212540 69080 212592 69086
rect 212540 69022 212592 69028
rect 212644 62830 212672 71862
rect 212632 62824 212684 62830
rect 212632 62766 212684 62772
rect 211252 10396 211304 10402
rect 211252 10338 211304 10344
rect 211172 6886 211752 6914
rect 210424 3460 210476 3466
rect 210424 3402 210476 3408
rect 210976 3392 211028 3398
rect 210976 3334 211028 3340
rect 209792 1958 209912 1986
rect 209792 480 209820 1958
rect 210988 480 211016 3334
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 6886
rect 213368 6248 213420 6254
rect 213368 6190 213420 6196
rect 213380 480 213408 6190
rect 213932 3534 213960 71878
rect 214116 71862 214190 71890
rect 214978 71936 215030 71942
rect 215818 71890 215846 72148
rect 214978 71878 215030 71884
rect 215312 71862 215846 71890
rect 216646 71890 216674 72148
rect 217474 71890 217502 72148
rect 218302 71890 218330 72148
rect 219130 71890 219158 72148
rect 219958 71890 219986 72148
rect 216646 71862 216720 71890
rect 214012 62824 214064 62830
rect 214012 62766 214064 62772
rect 214024 16574 214052 62766
rect 214116 57254 214144 71862
rect 214104 57248 214156 57254
rect 214104 57190 214156 57196
rect 214024 16546 214512 16574
rect 213920 3528 213972 3534
rect 213920 3470 213972 3476
rect 214484 480 214512 16546
rect 215312 6186 215340 71862
rect 216692 14482 216720 71862
rect 217428 71862 217502 71890
rect 218072 71862 218330 71890
rect 218532 71862 219158 71890
rect 219544 71862 219986 71890
rect 220786 71890 220814 72148
rect 221614 71890 221642 72148
rect 222442 71890 222470 72148
rect 223270 71890 223298 72148
rect 224098 71890 224126 72148
rect 220786 71862 220952 71890
rect 217324 70168 217376 70174
rect 217324 70110 217376 70116
rect 216680 14476 216732 14482
rect 216680 14418 216732 14424
rect 215300 6180 215352 6186
rect 215300 6122 215352 6128
rect 217336 4010 217364 70110
rect 217428 69766 217456 71862
rect 217416 69760 217468 69766
rect 217416 69702 217468 69708
rect 218072 11762 218100 71862
rect 218532 64874 218560 71862
rect 219440 69692 219492 69698
rect 219440 69634 219492 69640
rect 218164 64846 218560 64874
rect 218164 50386 218192 64846
rect 218152 50380 218204 50386
rect 218152 50322 218204 50328
rect 218152 49020 218204 49026
rect 218152 48962 218204 48968
rect 218060 11756 218112 11762
rect 218060 11698 218112 11704
rect 218164 6914 218192 48962
rect 218072 6886 218192 6914
rect 217324 4004 217376 4010
rect 217324 3946 217376 3952
rect 216864 3936 216916 3942
rect 216864 3878 216916 3884
rect 215668 3868 215720 3874
rect 215668 3810 215720 3816
rect 215680 480 215708 3810
rect 216876 480 216904 3878
rect 218072 480 218100 6886
rect 219256 3460 219308 3466
rect 219256 3402 219308 3408
rect 219268 480 219296 3402
rect 219452 490 219480 69634
rect 219544 3602 219572 71862
rect 220820 64388 220872 64394
rect 220820 64330 220872 64336
rect 220832 16574 220860 64330
rect 220924 64190 220952 71862
rect 221016 71862 221642 71890
rect 222396 71862 222470 71890
rect 223224 71862 223298 71890
rect 223592 71862 224126 71890
rect 224926 71890 224954 72148
rect 225754 71890 225782 72148
rect 226582 71890 226610 72148
rect 227410 71890 227438 72148
rect 228238 71890 228266 72148
rect 224926 71862 225000 71890
rect 221016 64258 221044 71862
rect 221464 70032 221516 70038
rect 221464 69974 221516 69980
rect 221004 64252 221056 64258
rect 221004 64194 221056 64200
rect 220912 64184 220964 64190
rect 220912 64126 220964 64132
rect 220832 16546 221136 16574
rect 219532 3596 219584 3602
rect 219532 3538 219584 3544
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 219452 462 220032 490
rect 220004 354 220032 462
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 221476 4078 221504 69974
rect 222396 69902 222424 71862
rect 222384 69896 222436 69902
rect 222384 69838 222436 69844
rect 223224 68406 223252 71862
rect 223212 68400 223264 68406
rect 223212 68342 223264 68348
rect 223592 4826 223620 71862
rect 224972 69086 225000 71862
rect 225708 71862 225782 71890
rect 226536 71862 226610 71890
rect 227364 71862 227438 71890
rect 228192 71862 228266 71890
rect 229066 71890 229094 72148
rect 229894 71890 229922 72148
rect 230722 71890 230750 72148
rect 231550 71890 231578 72148
rect 232378 71890 232406 72148
rect 229066 71862 229140 71890
rect 225604 69896 225656 69902
rect 225604 69838 225656 69844
rect 224224 69080 224276 69086
rect 224224 69022 224276 69028
rect 224960 69080 225012 69086
rect 224960 69022 225012 69028
rect 223672 44872 223724 44878
rect 223672 44814 223724 44820
rect 223580 4820 223632 4826
rect 223580 4762 223632 4768
rect 221464 4072 221516 4078
rect 221464 4014 221516 4020
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 222764 480 222792 3334
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223684 354 223712 44814
rect 224236 3670 224264 69022
rect 224960 65816 225012 65822
rect 224960 65758 225012 65764
rect 224972 16574 225000 65758
rect 224972 16546 225184 16574
rect 224224 3664 224276 3670
rect 224224 3606 224276 3612
rect 225156 480 225184 16546
rect 225616 3738 225644 69838
rect 225708 65686 225736 71862
rect 226536 69970 226564 71862
rect 227364 70106 227392 71862
rect 227352 70100 227404 70106
rect 227352 70042 227404 70048
rect 226524 69964 226576 69970
rect 226524 69906 226576 69912
rect 227720 68332 227772 68338
rect 227720 68274 227772 68280
rect 225696 65680 225748 65686
rect 225696 65622 225748 65628
rect 227732 16574 227760 68274
rect 228192 67046 228220 71862
rect 229112 70174 229140 71862
rect 229848 71862 229922 71890
rect 230492 71862 230750 71890
rect 230952 71862 231578 71890
rect 232332 71862 232406 71890
rect 233206 71890 233234 72148
rect 234034 71890 234062 72148
rect 234862 71890 234890 72148
rect 235690 71890 235718 72148
rect 236518 71890 236546 72148
rect 233206 71862 233280 71890
rect 229100 70168 229152 70174
rect 229100 70110 229152 70116
rect 228364 69964 228416 69970
rect 228364 69906 228416 69912
rect 228180 67040 228232 67046
rect 228180 66982 228232 66988
rect 227732 16546 228312 16574
rect 225604 3732 225656 3738
rect 225604 3674 225656 3680
rect 227536 3596 227588 3602
rect 227536 3538 227588 3544
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 226352 480 226380 3470
rect 227548 480 227576 3538
rect 223918 354 224030 480
rect 223684 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228376 3534 228404 69906
rect 229848 69902 229876 71862
rect 229836 69896 229888 69902
rect 229836 69838 229888 69844
rect 229100 69760 229152 69766
rect 229100 69702 229152 69708
rect 229112 16574 229140 69702
rect 229744 69080 229796 69086
rect 229744 69022 229796 69028
rect 229112 16546 229416 16574
rect 228364 3528 228416 3534
rect 228364 3470 228416 3476
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 229756 3806 229784 69022
rect 230492 7682 230520 71862
rect 230952 64874 230980 71862
rect 232332 69834 232360 71862
rect 232320 69828 232372 69834
rect 232320 69770 232372 69776
rect 233252 68474 233280 71862
rect 233988 71862 234062 71890
rect 234816 71862 234890 71890
rect 235644 71862 235718 71890
rect 236472 71862 236546 71890
rect 237346 71890 237374 72148
rect 238174 71890 238202 72148
rect 239002 71890 239030 72148
rect 239830 71890 239858 72148
rect 240658 71890 240686 72148
rect 237346 71862 237420 71890
rect 233332 70372 233384 70378
rect 233332 70314 233384 70320
rect 233240 68468 233292 68474
rect 233240 68410 233292 68416
rect 233344 64874 233372 70314
rect 233988 70038 234016 71862
rect 233976 70032 234028 70038
rect 233976 69974 234028 69980
rect 233884 69556 233936 69562
rect 233884 69498 233936 69504
rect 230584 64846 230980 64874
rect 233252 64846 233372 64874
rect 230584 13122 230612 64846
rect 231860 42084 231912 42090
rect 231860 42026 231912 42032
rect 230572 13116 230624 13122
rect 230572 13058 230624 13064
rect 230480 7676 230532 7682
rect 230480 7618 230532 7624
rect 229744 3800 229796 3806
rect 229744 3742 229796 3748
rect 231032 3664 231084 3670
rect 231032 3606 231084 3612
rect 231044 480 231072 3606
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 42026
rect 233252 16574 233280 64846
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 233896 3874 233924 69498
rect 234816 69086 234844 71862
rect 235264 69896 235316 69902
rect 235264 69838 235316 69844
rect 234804 69080 234856 69086
rect 234804 69022 234856 69028
rect 235276 3942 235304 69838
rect 235644 67114 235672 71862
rect 236000 69828 236052 69834
rect 236000 69770 236052 69776
rect 235632 67108 235684 67114
rect 235632 67050 235684 67056
rect 236012 16574 236040 69770
rect 236472 65550 236500 71862
rect 236460 65544 236512 65550
rect 236460 65486 236512 65492
rect 236012 16546 236592 16574
rect 235816 4820 235868 4826
rect 235816 4762 235868 4768
rect 235264 3936 235316 3942
rect 235264 3878 235316 3884
rect 233884 3868 233936 3874
rect 233884 3810 233936 3816
rect 234620 3732 234672 3738
rect 234620 3674 234672 3680
rect 234632 480 234660 3674
rect 235828 480 235856 4762
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237392 6254 237420 71862
rect 237484 71862 238202 71890
rect 238956 71862 239030 71890
rect 239784 71862 239858 71890
rect 240152 71862 240686 71890
rect 241486 71890 241514 72148
rect 242314 71890 242342 72148
rect 243142 71890 243170 72148
rect 243970 71890 243998 72148
rect 244798 71890 244826 72148
rect 241486 71862 241560 71890
rect 237484 62830 237512 71862
rect 238024 70236 238076 70242
rect 238024 70178 238076 70184
rect 237472 62824 237524 62830
rect 237472 62766 237524 62772
rect 237380 6248 237432 6254
rect 237380 6190 237432 6196
rect 238036 3466 238064 70178
rect 238956 69562 238984 71862
rect 239784 69902 239812 71862
rect 239772 69896 239824 69902
rect 239772 69838 239824 69844
rect 238944 69556 238996 69562
rect 238944 69498 238996 69504
rect 239404 69148 239456 69154
rect 239404 69090 239456 69096
rect 238760 66904 238812 66910
rect 238760 66846 238812 66852
rect 238772 16574 238800 66846
rect 238772 16546 239352 16574
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238024 3460 238076 3466
rect 238024 3402 238076 3408
rect 238128 480 238156 3742
rect 239324 480 239352 16546
rect 239416 3602 239444 69090
rect 240152 49026 240180 71862
rect 241532 70242 241560 71862
rect 242268 71862 242342 71890
rect 243004 71862 243170 71890
rect 243924 71862 243998 71890
rect 244292 71862 244826 71890
rect 245626 71890 245654 72148
rect 246454 71890 246482 72148
rect 247282 71890 247310 72148
rect 248110 71890 248138 72148
rect 248938 71890 248966 72148
rect 245626 71862 245700 71890
rect 241520 70236 241572 70242
rect 241520 70178 241572 70184
rect 242268 69698 242296 71862
rect 242256 69692 242308 69698
rect 242256 69634 242308 69640
rect 242900 69692 242952 69698
rect 242900 69634 242952 69640
rect 242256 69556 242308 69562
rect 242256 69498 242308 69504
rect 242164 69080 242216 69086
rect 242164 69022 242216 69028
rect 240140 49020 240192 49026
rect 240140 48962 240192 48968
rect 241704 4888 241756 4894
rect 241704 4830 241756 4836
rect 239404 3596 239456 3602
rect 239404 3538 239456 3544
rect 240508 3460 240560 3466
rect 240508 3402 240560 3408
rect 240520 480 240548 3402
rect 241716 480 241744 4830
rect 242176 3534 242204 69022
rect 242268 3670 242296 69498
rect 242912 11762 242940 69634
rect 243004 64394 243032 71862
rect 243924 69086 243952 71862
rect 243912 69080 243964 69086
rect 243912 69022 243964 69028
rect 242992 64388 243044 64394
rect 242992 64330 243044 64336
rect 242992 64184 243044 64190
rect 242992 64126 243044 64132
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 243004 6914 243032 64126
rect 244292 44878 244320 71862
rect 245672 65822 245700 71862
rect 246408 71862 246482 71890
rect 247236 71862 247310 71890
rect 248064 71862 248138 71890
rect 248892 71862 248966 71890
rect 249766 71890 249794 72148
rect 250594 71890 250622 72148
rect 251422 71890 251450 72148
rect 252250 71890 252278 72148
rect 253078 71890 253106 72148
rect 249766 71862 249840 71890
rect 246304 70304 246356 70310
rect 246304 70246 246356 70252
rect 245660 65816 245712 65822
rect 245660 65758 245712 65764
rect 245660 65544 245712 65550
rect 245660 65486 245712 65492
rect 244280 44872 244332 44878
rect 244280 44814 244332 44820
rect 245672 16574 245700 65486
rect 245672 16546 245976 16574
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242912 6886 243032 6914
rect 242256 3664 242308 3670
rect 242256 3606 242308 3612
rect 242164 3528 242216 3534
rect 242164 3470 242216 3476
rect 242912 480 242940 6886
rect 244108 480 244136 11698
rect 245200 3528 245252 3534
rect 245200 3470 245252 3476
rect 245212 480 245240 3470
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246316 3738 246344 70246
rect 246408 69970 246436 71862
rect 246396 69964 246448 69970
rect 246396 69906 246448 69912
rect 247040 69964 247092 69970
rect 247040 69906 247092 69912
rect 247052 16574 247080 69906
rect 247236 69154 247264 71862
rect 247684 70236 247736 70242
rect 247684 70178 247736 70184
rect 247224 69148 247276 69154
rect 247224 69090 247276 69096
rect 247052 16546 247632 16574
rect 246304 3732 246356 3738
rect 246304 3674 246356 3680
rect 247604 480 247632 16546
rect 247696 3806 247724 70178
rect 248064 68338 248092 71862
rect 248420 70032 248472 70038
rect 248420 69974 248472 69980
rect 248052 68332 248104 68338
rect 248052 68274 248104 68280
rect 247684 3800 247736 3806
rect 247684 3742 247736 3748
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 69974
rect 248892 69766 248920 71862
rect 248880 69760 248932 69766
rect 248880 69702 248932 69708
rect 249812 69562 249840 71862
rect 249904 71862 250622 71890
rect 251376 71862 251450 71890
rect 252204 71862 252278 71890
rect 252572 71862 253106 71890
rect 253906 71890 253934 72148
rect 254734 71890 254762 72148
rect 255562 71890 255590 72148
rect 256390 71890 256418 72148
rect 257218 71890 257246 72148
rect 253906 71862 253980 71890
rect 249800 69556 249852 69562
rect 249800 69498 249852 69504
rect 249800 68332 249852 68338
rect 249800 68274 249852 68280
rect 249812 16574 249840 68274
rect 249904 42090 249932 71862
rect 251376 70378 251404 71862
rect 251364 70372 251416 70378
rect 251364 70314 251416 70320
rect 252204 70310 252232 71862
rect 252192 70304 252244 70310
rect 252192 70246 252244 70252
rect 251272 69896 251324 69902
rect 251272 69838 251324 69844
rect 251180 69760 251232 69766
rect 251180 69702 251232 69708
rect 249892 42084 249944 42090
rect 249892 42026 249944 42032
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3602 251220 69702
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 251284 3482 251312 69838
rect 252572 4826 252600 71862
rect 253952 69834 253980 71862
rect 254688 71862 254762 71890
rect 255516 71862 255590 71890
rect 256344 71862 256418 71890
rect 256804 71862 257246 71890
rect 258046 71890 258074 72148
rect 258874 71890 258902 72148
rect 259702 71890 259730 72148
rect 260530 71890 260558 72148
rect 261358 71890 261386 72148
rect 258046 71862 258120 71890
rect 254688 70242 254716 71862
rect 254676 70236 254728 70242
rect 254676 70178 254728 70184
rect 254032 70100 254084 70106
rect 254032 70042 254084 70048
rect 253940 69828 253992 69834
rect 253940 69770 253992 69776
rect 253204 68468 253256 68474
rect 253204 68410 253256 68416
rect 252560 4820 252612 4826
rect 252560 4762 252612 4768
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253216 3466 253244 68410
rect 254044 64874 254072 70042
rect 255320 69828 255372 69834
rect 255320 69770 255372 69776
rect 253952 64846 254072 64874
rect 253952 16574 253980 64846
rect 255332 16574 255360 69770
rect 255516 66910 255544 71862
rect 256344 68474 256372 71862
rect 256700 70168 256752 70174
rect 256700 70110 256752 70116
rect 256332 68468 256384 68474
rect 256332 68410 256384 68416
rect 255504 66904 255556 66910
rect 255504 66846 255556 66852
rect 255964 66292 256016 66298
rect 255964 66234 256016 66240
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 253480 4820 253532 4826
rect 253480 4762 253532 4768
rect 253204 3460 253256 3466
rect 253204 3402 253256 3408
rect 253492 480 253520 4762
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 255976 3534 256004 66234
rect 255964 3528 256016 3534
rect 255964 3470 256016 3476
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 70110
rect 256804 4894 256832 71862
rect 258092 64190 258120 71862
rect 258828 71862 258902 71890
rect 259656 71862 259730 71890
rect 260484 71862 260558 71890
rect 261312 71862 261386 71890
rect 262186 71890 262214 72148
rect 263014 71890 263042 72148
rect 263842 71890 263870 72148
rect 264670 71890 264698 72148
rect 265498 71890 265526 72148
rect 262186 71862 262260 71890
rect 258828 69698 258856 71862
rect 258816 69692 258868 69698
rect 258816 69634 258868 69640
rect 259460 69692 259512 69698
rect 259460 69634 259512 69640
rect 258080 64184 258132 64190
rect 258080 64126 258132 64132
rect 259472 11762 259500 69634
rect 259656 66298 259684 71862
rect 259644 66292 259696 66298
rect 259644 66234 259696 66240
rect 259552 65680 259604 65686
rect 259552 65622 259604 65628
rect 259460 11756 259512 11762
rect 259460 11698 259512 11704
rect 259564 6914 259592 65622
rect 260484 65550 260512 71862
rect 260840 70236 260892 70242
rect 260840 70178 260892 70184
rect 260472 65544 260524 65550
rect 260472 65486 260524 65492
rect 260852 16574 260880 70178
rect 261312 69970 261340 71862
rect 262232 70038 262260 71862
rect 262968 71862 263042 71890
rect 263796 71862 263870 71890
rect 264624 71862 264698 71890
rect 265084 71862 265526 71890
rect 266326 71890 266354 72148
rect 267154 71890 267182 72148
rect 267982 71890 268010 72148
rect 268810 71890 268838 72148
rect 269638 71890 269666 72148
rect 266326 71862 266400 71890
rect 262220 70032 262272 70038
rect 262220 69974 262272 69980
rect 261300 69964 261352 69970
rect 261300 69906 261352 69912
rect 261484 69284 261536 69290
rect 261484 69226 261536 69232
rect 260852 16546 261432 16574
rect 260656 11756 260708 11762
rect 260656 11698 260708 11704
rect 259472 6886 259592 6914
rect 256792 4888 256844 4894
rect 256792 4830 256844 4836
rect 258264 3596 258316 3602
rect 258264 3538 258316 3544
rect 258276 480 258304 3538
rect 259472 480 259500 6886
rect 260668 480 260696 11698
rect 261404 3482 261432 16546
rect 261496 3602 261524 69226
rect 262968 68338 262996 71862
rect 263600 70032 263652 70038
rect 263600 69974 263652 69980
rect 262956 68332 263008 68338
rect 262956 68274 263008 68280
rect 263612 16574 263640 69974
rect 263796 69902 263824 71862
rect 263784 69896 263836 69902
rect 263784 69838 263836 69844
rect 264624 69766 264652 71862
rect 264980 69896 265032 69902
rect 264980 69838 265032 69844
rect 264612 69760 264664 69766
rect 264612 69702 264664 69708
rect 263612 16546 264192 16574
rect 262956 4140 263008 4146
rect 262956 4082 263008 4088
rect 261484 3596 261536 3602
rect 261484 3538 261536 3544
rect 261404 3454 261800 3482
rect 261772 480 261800 3454
rect 262968 480 262996 4082
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 69838
rect 265084 4826 265112 71862
rect 266372 70106 266400 71862
rect 267108 71862 267182 71890
rect 267936 71862 268010 71890
rect 268764 71862 268838 71890
rect 269592 71862 269666 71890
rect 270466 71890 270494 72148
rect 271294 71890 271322 72148
rect 272122 71890 272150 72148
rect 272950 71890 272978 72148
rect 273778 71890 273806 72148
rect 270466 71862 270540 71890
rect 266360 70100 266412 70106
rect 266360 70042 266412 70048
rect 266360 69964 266412 69970
rect 266360 69906 266412 69912
rect 266372 16574 266400 69906
rect 267108 69834 267136 71862
rect 267936 70174 267964 71862
rect 267924 70168 267976 70174
rect 267924 70110 267976 70116
rect 267096 69828 267148 69834
rect 267096 69770 267148 69776
rect 267740 69352 267792 69358
rect 267740 69294 267792 69300
rect 266372 16546 266584 16574
rect 265072 4820 265124 4826
rect 265072 4762 265124 4768
rect 266556 480 266584 16546
rect 267752 3602 267780 69294
rect 268764 69290 268792 71862
rect 268752 69284 268804 69290
rect 268752 69226 268804 69232
rect 267832 69216 267884 69222
rect 267832 69158 267884 69164
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 267844 3482 267872 69158
rect 269120 69148 269172 69154
rect 269120 69090 269172 69096
rect 269132 16574 269160 69090
rect 269592 65686 269620 71862
rect 270512 69698 270540 71862
rect 271248 71862 271322 71890
rect 272076 71862 272150 71890
rect 272904 71862 272978 71890
rect 273732 71862 273806 71890
rect 274606 71890 274634 72148
rect 275434 71890 275462 72148
rect 276262 71890 276290 72148
rect 277090 71890 277118 72148
rect 277918 71890 277946 72148
rect 274606 71862 274680 71890
rect 271248 70242 271276 71862
rect 271236 70236 271288 70242
rect 271236 70178 271288 70184
rect 270500 69692 270552 69698
rect 270500 69634 270552 69640
rect 270500 69556 270552 69562
rect 270500 69498 270552 69504
rect 269764 69080 269816 69086
rect 269764 69022 269816 69028
rect 269580 65680 269632 65686
rect 269580 65622 269632 65628
rect 269132 16546 269712 16574
rect 268476 3596 268528 3602
rect 268476 3538 268528 3544
rect 267752 3454 267872 3482
rect 267752 480 267780 3454
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3538
rect 269684 3482 269712 16546
rect 269776 4146 269804 69022
rect 270512 16574 270540 69498
rect 272076 69086 272104 71862
rect 272904 70038 272932 71862
rect 272892 70032 272944 70038
rect 272892 69974 272944 69980
rect 273260 70032 273312 70038
rect 273260 69974 273312 69980
rect 272064 69080 272116 69086
rect 272064 69022 272116 69028
rect 270512 16546 270816 16574
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 269684 3454 270080 3482
rect 270052 480 270080 3454
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 272444 480 272472 3470
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 69974
rect 273732 69902 273760 71862
rect 274652 69970 274680 71862
rect 275388 71862 275462 71890
rect 276216 71862 276290 71890
rect 277044 71862 277118 71890
rect 277872 71862 277946 71890
rect 278746 71890 278774 72148
rect 279574 71890 279602 72148
rect 280402 71890 280430 72148
rect 281230 71890 281258 72148
rect 282058 71890 282086 72148
rect 278746 71862 278820 71890
rect 274640 69964 274692 69970
rect 274640 69906 274692 69912
rect 273720 69896 273772 69902
rect 273720 69838 273772 69844
rect 273904 69896 273956 69902
rect 273904 69838 273956 69844
rect 273916 3534 273944 69838
rect 274640 69692 274692 69698
rect 274640 69634 274692 69640
rect 274652 16574 274680 69634
rect 275388 69222 275416 71862
rect 276216 69358 276244 71862
rect 276204 69352 276256 69358
rect 276204 69294 276256 69300
rect 275376 69216 275428 69222
rect 275376 69158 275428 69164
rect 277044 69154 277072 71862
rect 277872 69562 277900 71862
rect 278792 69902 278820 71862
rect 279528 71862 279602 71890
rect 280356 71862 280430 71890
rect 281184 71862 281258 71890
rect 282012 71862 282086 71890
rect 282886 71890 282914 72148
rect 283714 71890 283742 72148
rect 284542 71890 284570 72148
rect 285370 71890 285398 72148
rect 286198 71890 286226 72148
rect 282886 71862 282960 71890
rect 279528 70038 279556 71862
rect 279516 70032 279568 70038
rect 279516 69974 279568 69980
rect 278780 69896 278832 69902
rect 278780 69838 278832 69844
rect 280356 69698 280384 71862
rect 280344 69692 280396 69698
rect 280344 69634 280396 69640
rect 277860 69556 277912 69562
rect 277860 69498 277912 69504
rect 277400 69284 277452 69290
rect 277400 69226 277452 69232
rect 277032 69148 277084 69154
rect 277032 69090 277084 69096
rect 277412 16574 277440 69226
rect 280160 69216 280212 69222
rect 280160 69158 280212 69164
rect 278044 69148 278096 69154
rect 278044 69090 278096 69096
rect 274652 16546 274864 16574
rect 277412 16546 277992 16574
rect 273904 3528 273956 3534
rect 273904 3470 273956 3476
rect 274836 480 274864 16546
rect 276020 3868 276072 3874
rect 276020 3810 276072 3816
rect 276032 480 276060 3810
rect 277124 3732 277176 3738
rect 277124 3674 277176 3680
rect 277136 480 277164 3674
rect 277964 3482 277992 16546
rect 278056 3874 278084 69090
rect 279424 69080 279476 69086
rect 279424 69022 279476 69028
rect 278044 3868 278096 3874
rect 278044 3810 278096 3816
rect 279436 3738 279464 69022
rect 280172 16574 280200 69158
rect 281184 69154 281212 71862
rect 281172 69148 281224 69154
rect 281172 69090 281224 69096
rect 281540 69148 281592 69154
rect 281540 69090 281592 69096
rect 280172 16546 280752 16574
rect 279424 3732 279476 3738
rect 279424 3674 279476 3680
rect 279516 3732 279568 3738
rect 279516 3674 279568 3680
rect 277964 3454 278360 3482
rect 278332 480 278360 3454
rect 279528 480 279556 3674
rect 280724 480 280752 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 354 281580 69090
rect 282012 69086 282040 71862
rect 282932 69290 282960 71862
rect 283116 71862 283742 71890
rect 284496 71862 284570 71890
rect 285324 71862 285398 71890
rect 285784 71862 286226 71890
rect 287026 71890 287054 72148
rect 287854 71890 287882 72148
rect 288682 71890 288710 72148
rect 289510 71890 289538 72148
rect 290338 71890 290366 72148
rect 287026 71862 287192 71890
rect 282920 69284 282972 69290
rect 282920 69226 282972 69232
rect 282000 69080 282052 69086
rect 282000 69022 282052 69028
rect 283116 3738 283144 71862
rect 284300 69284 284352 69290
rect 284300 69226 284352 69232
rect 284312 16574 284340 69226
rect 284496 69222 284524 71862
rect 284484 69216 284536 69222
rect 284484 69158 284536 69164
rect 285324 69154 285352 71862
rect 285680 69828 285732 69834
rect 285680 69770 285732 69776
rect 285312 69148 285364 69154
rect 285312 69090 285364 69096
rect 284312 16546 284984 16574
rect 284300 4140 284352 4146
rect 284300 4082 284352 4088
rect 283104 3732 283156 3738
rect 283104 3674 283156 3680
rect 283104 3596 283156 3602
rect 283104 3538 283156 3544
rect 283116 480 283144 3538
rect 284312 480 284340 4082
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 285692 3482 285720 69770
rect 285784 3602 285812 71862
rect 287060 69148 287112 69154
rect 287060 69090 287112 69096
rect 285772 3596 285824 3602
rect 285772 3538 285824 3544
rect 285692 3454 286640 3482
rect 286612 480 286640 3454
rect 287072 490 287100 69090
rect 287164 4146 287192 71862
rect 287808 71862 287882 71890
rect 288636 71862 288710 71890
rect 289464 71862 289538 71890
rect 290292 71862 290366 71890
rect 291166 71890 291194 72148
rect 291994 71890 292022 72148
rect 292822 71890 292850 72148
rect 293650 71890 293678 72148
rect 294478 71890 294506 72148
rect 291166 71862 291240 71890
rect 287808 69290 287836 71862
rect 288636 69834 288664 71862
rect 288624 69828 288676 69834
rect 288624 69770 288676 69776
rect 287796 69284 287848 69290
rect 287796 69226 287848 69232
rect 289464 69154 289492 71862
rect 289452 69148 289504 69154
rect 289452 69090 289504 69096
rect 290292 69086 290320 71862
rect 288440 69080 288492 69086
rect 288440 69022 288492 69028
rect 290280 69080 290332 69086
rect 290280 69022 290332 69028
rect 288452 16574 288480 69022
rect 288452 16546 289032 16574
rect 287152 4140 287204 4146
rect 287152 4082 287204 4088
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287072 462 287376 490
rect 289004 480 289032 16546
rect 291212 3466 291240 71862
rect 291396 71862 292022 71890
rect 292592 71862 292850 71890
rect 293144 71862 293678 71890
rect 293972 71862 294506 71890
rect 295306 71890 295334 72148
rect 296134 71890 296162 72148
rect 295306 71862 295380 71890
rect 290188 3460 290240 3466
rect 290188 3402 290240 3408
rect 291200 3460 291252 3466
rect 291200 3402 291252 3408
rect 290200 480 290228 3402
rect 291396 480 291424 71862
rect 292592 480 292620 71862
rect 293144 64874 293172 71862
rect 292684 64846 293172 64874
rect 292684 16574 292712 64846
rect 293972 16574 294000 71862
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 287348 354 287376 462
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295352 490 295380 71862
rect 295444 71862 296162 71890
rect 296812 71936 296864 71942
rect 296962 71890 296990 72148
rect 297790 71942 297818 72148
rect 296812 71878 296864 71884
rect 295444 3058 295472 71862
rect 296824 3466 296852 71878
rect 296916 71862 296990 71890
rect 297778 71936 297830 71942
rect 297778 71878 297830 71884
rect 298618 71890 298646 72148
rect 299446 71890 299474 72148
rect 300274 71890 300302 72148
rect 301102 72026 301130 72148
rect 300872 71998 301130 72026
rect 298618 71862 298692 71890
rect 299446 71862 299520 71890
rect 300274 71862 300348 71890
rect 296812 3460 296864 3466
rect 296812 3402 296864 3408
rect 295432 3052 295484 3058
rect 295432 2994 295484 3000
rect 296916 2990 296944 71862
rect 298664 69086 298692 71862
rect 299492 69154 299520 71862
rect 299480 69148 299532 69154
rect 299480 69090 299532 69096
rect 300320 69086 300348 71862
rect 300872 69290 300900 71998
rect 301930 71890 301958 72148
rect 302758 71890 302786 72148
rect 300964 71862 301958 71890
rect 302344 71862 302786 71890
rect 303586 71890 303614 72148
rect 304414 71890 304442 72148
rect 305242 71890 305270 72148
rect 303586 71862 303752 71890
rect 304414 71862 304488 71890
rect 300860 69284 300912 69290
rect 300860 69226 300912 69232
rect 300860 69148 300912 69154
rect 300860 69090 300912 69096
rect 298652 69080 298704 69086
rect 298652 69022 298704 69028
rect 299756 69080 299808 69086
rect 299756 69022 299808 69028
rect 300308 69080 300360 69086
rect 300308 69022 300360 69028
rect 299768 16574 299796 69022
rect 299768 16546 300808 16574
rect 299664 3460 299716 3466
rect 299664 3402 299716 3408
rect 297272 3052 297324 3058
rect 297272 2994 297324 3000
rect 296904 2984 296956 2990
rect 296904 2926 296956 2932
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295352 462 295656 490
rect 297284 480 297312 2994
rect 298468 2984 298520 2990
rect 298468 2926 298520 2932
rect 298480 480 298508 2926
rect 299676 480 299704 3402
rect 300780 480 300808 16546
rect 300872 2530 300900 69090
rect 300964 3534 300992 71862
rect 302240 69080 302292 69086
rect 302240 69022 302292 69028
rect 300952 3528 301004 3534
rect 300952 3470 301004 3476
rect 302252 3482 302280 69022
rect 302344 4146 302372 71862
rect 303620 69284 303672 69290
rect 303620 69226 303672 69232
rect 302332 4140 302384 4146
rect 302332 4082 302384 4088
rect 303528 4140 303580 4146
rect 303528 4082 303580 4088
rect 302252 3454 303200 3482
rect 300872 2502 301544 2530
rect 295628 354 295656 462
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 2502
rect 303172 480 303200 3454
rect 303540 3058 303568 4082
rect 303528 3052 303580 3058
rect 303528 2994 303580 3000
rect 303632 490 303660 69226
rect 303724 3738 303752 71862
rect 304460 69086 304488 71862
rect 305012 71862 305270 71890
rect 306070 71890 306098 72148
rect 306898 71890 306926 72148
rect 306070 71862 306144 71890
rect 304448 69080 304500 69086
rect 304448 69022 304500 69028
rect 303712 3732 303764 3738
rect 303712 3674 303764 3680
rect 305012 3670 305040 71862
rect 306116 69902 306144 71862
rect 306484 71862 306926 71890
rect 307726 71890 307754 72148
rect 308554 71890 308582 72148
rect 309140 71936 309192 71942
rect 307726 71862 307800 71890
rect 308554 71862 308628 71890
rect 309382 71890 309410 72148
rect 310210 71942 310238 72148
rect 309140 71878 309192 71884
rect 306104 69896 306156 69902
rect 306104 69838 306156 69844
rect 305644 69080 305696 69086
rect 305644 69022 305696 69028
rect 305656 3942 305684 69022
rect 305644 3936 305696 3942
rect 305644 3878 305696 3884
rect 305000 3664 305052 3670
rect 305000 3606 305052 3612
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303632 462 303936 490
rect 305564 480 305592 3470
rect 306484 2990 306512 71862
rect 307024 69896 307076 69902
rect 307024 69838 307076 69844
rect 307036 3466 307064 69838
rect 307772 69086 307800 71862
rect 308600 69154 308628 71862
rect 308588 69148 308640 69154
rect 308588 69090 308640 69096
rect 307760 69080 307812 69086
rect 307760 69022 307812 69028
rect 309048 3936 309100 3942
rect 309048 3878 309100 3884
rect 307944 3732 307996 3738
rect 307944 3674 307996 3680
rect 307024 3460 307076 3466
rect 307024 3402 307076 3408
rect 306748 3052 306800 3058
rect 306748 2994 306800 3000
rect 306472 2984 306524 2990
rect 306472 2926 306524 2932
rect 306760 480 306788 2994
rect 307956 480 307984 3674
rect 309060 480 309088 3878
rect 309152 3126 309180 71878
rect 309336 71862 309410 71890
rect 310198 71936 310250 71942
rect 311038 71890 311066 72148
rect 310198 71878 310250 71884
rect 310532 71862 311066 71890
rect 311866 71890 311894 72148
rect 312694 71890 312722 72148
rect 313522 71890 313550 72148
rect 314350 71890 314378 72148
rect 315178 71890 315206 72148
rect 311866 71862 311940 71890
rect 312694 71862 312768 71890
rect 309336 3262 309364 71862
rect 309784 69080 309836 69086
rect 309784 69022 309836 69028
rect 309796 3534 309824 69022
rect 310244 3664 310296 3670
rect 310244 3606 310296 3612
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 309324 3256 309376 3262
rect 309324 3198 309376 3204
rect 309140 3120 309192 3126
rect 309140 3062 309192 3068
rect 310256 480 310284 3606
rect 310532 3398 310560 71862
rect 311912 69698 311940 71862
rect 311900 69692 311952 69698
rect 311900 69634 311952 69640
rect 311164 69148 311216 69154
rect 311164 69090 311216 69096
rect 310520 3392 310572 3398
rect 310520 3334 310572 3340
rect 311176 3330 311204 69090
rect 312740 69086 312768 71862
rect 313384 71862 313550 71890
rect 313660 71862 314378 71890
rect 314672 71862 315206 71890
rect 316006 71890 316034 72148
rect 316834 71890 316862 72148
rect 316006 71862 316080 71890
rect 312728 69080 312780 69086
rect 312728 69022 312780 69028
rect 313384 3466 313412 71862
rect 313660 3670 313688 71862
rect 313924 69080 313976 69086
rect 313924 69022 313976 69028
rect 313936 3942 313964 69022
rect 314672 4962 314700 71862
rect 316052 69086 316080 71862
rect 316144 71862 316862 71890
rect 317662 71890 317690 72148
rect 318490 71890 318518 72148
rect 319318 71890 319346 72148
rect 317662 71862 317736 71890
rect 316040 69080 316092 69086
rect 316040 69022 316092 69028
rect 314660 4956 314712 4962
rect 314660 4898 314712 4904
rect 313924 3936 313976 3942
rect 313924 3878 313976 3884
rect 316144 3874 316172 71862
rect 317708 69154 317736 71862
rect 317800 71862 318518 71890
rect 318904 71862 319346 71890
rect 320146 71890 320174 72148
rect 320974 71890 321002 72148
rect 321802 71890 321830 72148
rect 322630 71890 322658 72148
rect 323458 71890 323486 72148
rect 320146 71862 320220 71890
rect 317696 69148 317748 69154
rect 317696 69090 317748 69096
rect 316132 3868 316184 3874
rect 316132 3810 316184 3816
rect 313648 3664 313700 3670
rect 313648 3606 313700 3612
rect 317800 3602 317828 71862
rect 318800 69692 318852 69698
rect 318800 69634 318852 69640
rect 318064 69080 318116 69086
rect 318064 69022 318116 69028
rect 317788 3596 317840 3602
rect 317788 3538 317840 3544
rect 313832 3528 313884 3534
rect 313832 3470 313884 3476
rect 311440 3460 311492 3466
rect 311440 3402 311492 3408
rect 313372 3460 313424 3466
rect 313372 3402 313424 3408
rect 311164 3324 311216 3330
rect 311164 3266 311216 3272
rect 311452 480 311480 3402
rect 312636 2984 312688 2990
rect 312636 2926 312688 2932
rect 312648 480 312676 2926
rect 313844 480 313872 3470
rect 318076 3330 318104 69022
rect 318812 3482 318840 69634
rect 318904 3806 318932 71862
rect 320192 69970 320220 71862
rect 320284 71862 321002 71890
rect 321572 71862 321830 71890
rect 322032 71862 322658 71890
rect 323044 71862 323486 71890
rect 324286 71890 324314 72148
rect 325114 71890 325142 72148
rect 324286 71862 324636 71890
rect 320180 69964 320232 69970
rect 320180 69906 320232 69912
rect 318892 3800 318944 3806
rect 318892 3742 318944 3748
rect 320284 3738 320312 71862
rect 321572 3942 321600 71862
rect 322032 64874 322060 71862
rect 321664 64846 322060 64874
rect 321664 7750 321692 64846
rect 321652 7744 321704 7750
rect 321652 7686 321704 7692
rect 320916 3936 320968 3942
rect 320916 3878 320968 3884
rect 321560 3936 321612 3942
rect 321560 3878 321612 3884
rect 320272 3732 320324 3738
rect 320272 3674 320324 3680
rect 318812 3454 319760 3482
rect 318524 3392 318576 3398
rect 318524 3334 318576 3340
rect 315028 3324 315080 3330
rect 315028 3266 315080 3272
rect 318064 3324 318116 3330
rect 318064 3266 318116 3272
rect 315040 480 315068 3266
rect 316224 3256 316276 3262
rect 316224 3198 316276 3204
rect 316236 480 316264 3198
rect 317328 3120 317380 3126
rect 317328 3062 317380 3068
rect 317340 480 317368 3062
rect 318536 480 318564 3334
rect 319732 480 319760 3454
rect 320928 480 320956 3878
rect 323044 3534 323072 71862
rect 323584 69148 323636 69154
rect 323584 69090 323636 69096
rect 323596 4418 323624 69090
rect 324412 66224 324464 66230
rect 324412 66166 324464 66172
rect 324320 4956 324372 4962
rect 324320 4898 324372 4904
rect 323584 4412 323636 4418
rect 323584 4354 323636 4360
rect 323308 3664 323360 3670
rect 323308 3606 323360 3612
rect 323032 3528 323084 3534
rect 323032 3470 323084 3476
rect 322112 3460 322164 3466
rect 322112 3402 322164 3408
rect 322124 480 322152 3402
rect 323320 480 323348 3606
rect 324332 2530 324360 4898
rect 324424 4826 324452 66166
rect 324412 4820 324464 4826
rect 324412 4762 324464 4768
rect 324608 3670 324636 71862
rect 325068 71862 325142 71890
rect 325942 71890 325970 72148
rect 326770 71890 326798 72148
rect 327598 71890 327626 72148
rect 325942 71862 326016 71890
rect 325068 66230 325096 71862
rect 325988 69698 326016 71862
rect 326080 71862 326798 71890
rect 327092 71862 327626 71890
rect 328426 71890 328454 72148
rect 329254 71890 329282 72148
rect 330082 71890 330110 72148
rect 328426 71862 328500 71890
rect 325976 69692 326028 69698
rect 325976 69634 326028 69640
rect 325056 66224 325108 66230
rect 325056 66166 325108 66172
rect 324596 3664 324648 3670
rect 324596 3606 324648 3612
rect 326080 3466 326108 71862
rect 327092 6186 327120 71862
rect 327724 69964 327776 69970
rect 327724 69906 327776 69912
rect 327080 6180 327132 6186
rect 327080 6122 327132 6128
rect 327736 4214 327764 69906
rect 328472 9042 328500 71862
rect 328564 71862 329282 71890
rect 329852 71862 330110 71890
rect 330910 71890 330938 72148
rect 331738 71890 331766 72148
rect 330910 71862 330984 71890
rect 328460 9036 328512 9042
rect 328460 8978 328512 8984
rect 328000 4412 328052 4418
rect 328000 4354 328052 4360
rect 327724 4208 327776 4214
rect 327724 4150 327776 4156
rect 326804 3868 326856 3874
rect 326804 3810 326856 3816
rect 326068 3460 326120 3466
rect 326068 3402 326120 3408
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 324332 2502 324452 2530
rect 324424 480 324452 2502
rect 325620 480 325648 3266
rect 326816 480 326844 3810
rect 328012 480 328040 4354
rect 328564 3874 328592 71862
rect 329852 15910 329880 71862
rect 330956 69086 330984 71862
rect 331324 71862 331766 71890
rect 332566 71890 332594 72148
rect 333394 71890 333422 72148
rect 332566 71862 332640 71890
rect 330944 69080 330996 69086
rect 330944 69022 330996 69028
rect 329840 15904 329892 15910
rect 329840 15846 329892 15852
rect 328552 3868 328604 3874
rect 328552 3810 328604 3816
rect 330392 3800 330444 3806
rect 330392 3742 330444 3748
rect 329196 3596 329248 3602
rect 329196 3538 329248 3544
rect 329208 480 329236 3538
rect 330404 480 330432 3742
rect 331324 3602 331352 71862
rect 331864 69080 331916 69086
rect 331864 69022 331916 69028
rect 331876 7682 331904 69022
rect 331864 7676 331916 7682
rect 331864 7618 331916 7624
rect 332612 4894 332640 71862
rect 332704 71862 333422 71890
rect 334222 71890 334250 72148
rect 335050 71890 335078 72148
rect 334222 71862 334296 71890
rect 332704 10402 332732 71862
rect 334268 69902 334296 71862
rect 334360 71862 335078 71890
rect 335878 71890 335906 72148
rect 336706 71890 336734 72148
rect 337534 71890 337562 72148
rect 338362 71890 338390 72148
rect 339190 71890 339218 72148
rect 340018 71890 340046 72148
rect 335878 71862 335952 71890
rect 336706 71862 336780 71890
rect 334256 69896 334308 69902
rect 334256 69838 334308 69844
rect 332692 10396 332744 10402
rect 332692 10338 332744 10344
rect 334360 7614 334388 71862
rect 335924 69766 335952 71862
rect 336004 69896 336056 69902
rect 336004 69838 336056 69844
rect 335912 69760 335964 69766
rect 335912 69702 335964 69708
rect 335084 7744 335136 7750
rect 335084 7686 335136 7692
rect 334348 7608 334400 7614
rect 334348 7550 334400 7556
rect 332600 4888 332652 4894
rect 332600 4830 332652 4836
rect 331588 4208 331640 4214
rect 331588 4150 331640 4156
rect 331312 3596 331364 3602
rect 331312 3538 331364 3544
rect 331600 480 331628 4150
rect 333888 3936 333940 3942
rect 333888 3878 333940 3884
rect 332692 3732 332744 3738
rect 332692 3674 332744 3680
rect 332704 480 332732 3674
rect 333900 480 333928 3878
rect 335096 480 335124 7686
rect 336016 3942 336044 69838
rect 336096 69692 336148 69698
rect 336096 69634 336148 69640
rect 336108 5574 336136 69634
rect 336096 5568 336148 5574
rect 336096 5510 336148 5516
rect 336004 3936 336056 3942
rect 336004 3878 336056 3884
rect 336752 3806 336780 71862
rect 336844 71862 337562 71890
rect 338132 71862 338390 71890
rect 338500 71862 339218 71890
rect 339604 71862 340046 71890
rect 340846 71890 340874 72148
rect 341674 71890 341702 72148
rect 342502 71890 342530 72148
rect 343330 71890 343358 72148
rect 340846 71862 340920 71890
rect 336844 8974 336872 71862
rect 338132 11898 338160 71862
rect 338120 11892 338172 11898
rect 338120 11834 338172 11840
rect 336832 8968 336884 8974
rect 336832 8910 336884 8916
rect 336740 3800 336792 3806
rect 336740 3742 336792 3748
rect 338500 3670 338528 71862
rect 339604 4826 339632 71862
rect 339868 5568 339920 5574
rect 339868 5510 339920 5516
rect 338672 4820 338724 4826
rect 338672 4762 338724 4768
rect 339592 4820 339644 4826
rect 339592 4762 339644 4768
rect 337476 3664 337528 3670
rect 337476 3606 337528 3612
rect 338488 3664 338540 3670
rect 338488 3606 338540 3612
rect 336280 3528 336332 3534
rect 336280 3470 336332 3476
rect 336292 480 336320 3470
rect 337488 480 337516 3606
rect 338684 480 338712 4762
rect 339880 480 339908 5510
rect 340892 3738 340920 71862
rect 340984 71862 341702 71890
rect 342272 71862 342530 71890
rect 342640 71862 343358 71890
rect 344158 71890 344186 72148
rect 344986 71890 345014 72148
rect 345814 71890 345842 72148
rect 344158 71862 344232 71890
rect 344986 71862 345060 71890
rect 340984 16574 341012 71862
rect 340984 16546 341104 16574
rect 340880 3732 340932 3738
rect 340880 3674 340932 3680
rect 341076 3534 341104 16546
rect 342272 10334 342300 71862
rect 342640 64874 342668 71862
rect 344204 69698 344232 71862
rect 344192 69692 344244 69698
rect 344192 69634 344244 69640
rect 345032 69154 345060 71862
rect 345124 71862 345842 71890
rect 346492 71936 346544 71942
rect 346642 71890 346670 72148
rect 347470 71942 347498 72148
rect 346492 71878 346544 71884
rect 345020 69148 345072 69154
rect 345020 69090 345072 69096
rect 342364 64846 342668 64874
rect 342364 11830 342392 64846
rect 345124 14482 345152 71862
rect 345664 69760 345716 69766
rect 345664 69702 345716 69708
rect 345296 15904 345348 15910
rect 345296 15846 345348 15852
rect 345112 14476 345164 14482
rect 345112 14418 345164 14424
rect 342352 11824 342404 11830
rect 342352 11766 342404 11772
rect 342260 10328 342312 10334
rect 342260 10270 342312 10276
rect 343364 9036 343416 9042
rect 343364 8978 343416 8984
rect 342168 6180 342220 6186
rect 342168 6122 342220 6128
rect 341064 3528 341116 3534
rect 341064 3470 341116 3476
rect 340972 3460 341024 3466
rect 340972 3402 341024 3408
rect 340984 480 341012 3402
rect 342180 480 342208 6122
rect 343376 480 343404 8978
rect 344560 3868 344612 3874
rect 344560 3810 344612 3816
rect 344572 480 344600 3810
rect 303908 354 303936 462
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 15846
rect 345676 13054 345704 69702
rect 345664 13048 345716 13054
rect 345664 12990 345716 12996
rect 346504 6458 346532 71878
rect 346596 71862 346670 71890
rect 347458 71936 347510 71942
rect 347458 71878 347510 71884
rect 348298 71890 348326 72148
rect 349126 71890 349154 72148
rect 349954 71890 349982 72148
rect 348298 71862 348372 71890
rect 349126 71862 349200 71890
rect 346492 6452 346544 6458
rect 346492 6394 346544 6400
rect 346596 3398 346624 71862
rect 348344 69086 348372 71862
rect 349172 69766 349200 71862
rect 349264 71862 349982 71890
rect 350782 71890 350810 72148
rect 351610 71890 351638 72148
rect 352438 71890 352466 72148
rect 350782 71862 350856 71890
rect 349160 69760 349212 69766
rect 349160 69702 349212 69708
rect 348332 69080 348384 69086
rect 348332 69022 348384 69028
rect 349160 10396 349212 10402
rect 349160 10338 349212 10344
rect 346952 7676 347004 7682
rect 346952 7618 347004 7624
rect 346584 3392 346636 3398
rect 346584 3334 346636 3340
rect 346964 480 346992 7618
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 348068 480 348096 3538
rect 349172 3466 349200 10338
rect 349264 6186 349292 71862
rect 350828 69902 350856 71862
rect 350920 71862 351638 71890
rect 351932 71862 352466 71890
rect 353266 71890 353294 72148
rect 354094 71890 354122 72148
rect 354922 71890 354950 72148
rect 353266 71862 353340 71890
rect 354094 71862 354168 71890
rect 350816 69896 350868 69902
rect 350816 69838 350868 69844
rect 349804 69148 349856 69154
rect 349804 69090 349856 69096
rect 349252 6180 349304 6186
rect 349252 6122 349304 6128
rect 349816 4962 349844 69090
rect 349804 4956 349856 4962
rect 349804 4898 349856 4904
rect 349252 4888 349304 4894
rect 349252 4830 349304 4836
rect 349160 3460 349212 3466
rect 349160 3402 349212 3408
rect 349264 480 349292 4830
rect 350920 3602 350948 71862
rect 351184 69080 351236 69086
rect 351184 69022 351236 69028
rect 351196 13394 351224 69022
rect 351184 13388 351236 13394
rect 351184 13330 351236 13336
rect 351932 7818 351960 71862
rect 353312 15910 353340 71862
rect 354140 69834 354168 71862
rect 354692 71862 354950 71890
rect 355750 71890 355778 72148
rect 356578 71890 356606 72148
rect 357406 71890 357434 72148
rect 358234 71890 358262 72148
rect 359062 72026 359090 72148
rect 359062 71998 359136 72026
rect 355750 71862 355824 71890
rect 356578 71862 356652 71890
rect 357406 71862 357480 71890
rect 358234 71862 358308 71890
rect 354128 69828 354180 69834
rect 354128 69770 354180 69776
rect 353300 15904 353352 15910
rect 353300 15846 353352 15852
rect 353576 13048 353628 13054
rect 353576 12990 353628 12996
rect 351920 7812 351972 7818
rect 351920 7754 351972 7760
rect 352840 7608 352892 7614
rect 352840 7550 352892 7556
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 350908 3596 350960 3602
rect 350908 3538 350960 3544
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 350460 480 350488 3402
rect 351656 480 351684 3878
rect 352852 480 352880 7550
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 12990
rect 354692 7750 354720 71862
rect 355324 69896 355376 69902
rect 355324 69838 355376 69844
rect 354680 7744 354732 7750
rect 354680 7686 354732 7692
rect 355336 4894 355364 69838
rect 355796 69086 355824 71862
rect 356624 69154 356652 71862
rect 356612 69148 356664 69154
rect 356612 69090 356664 69096
rect 357452 69086 357480 71862
rect 358280 69698 358308 71862
rect 359108 70106 359136 71998
rect 359890 71890 359918 72148
rect 360718 71890 360746 72148
rect 359292 71862 359918 71890
rect 360212 71862 360746 71890
rect 361546 71890 361574 72148
rect 362374 71890 362402 72148
rect 363202 71890 363230 72148
rect 361546 71862 361620 71890
rect 362374 71862 362448 71890
rect 359096 70100 359148 70106
rect 359096 70042 359148 70048
rect 358084 69692 358136 69698
rect 358084 69634 358136 69640
rect 358268 69692 358320 69698
rect 358268 69634 358320 69640
rect 355784 69080 355836 69086
rect 355784 69022 355836 69028
rect 356704 69080 356756 69086
rect 356704 69022 356756 69028
rect 357440 69080 357492 69086
rect 357440 69022 357492 69028
rect 356716 11762 356744 69022
rect 357532 11892 357584 11898
rect 357532 11834 357584 11840
rect 356704 11756 356756 11762
rect 356704 11698 356756 11704
rect 356336 8968 356388 8974
rect 356336 8910 356388 8916
rect 355324 4888 355376 4894
rect 355324 4830 355376 4836
rect 355232 3800 355284 3806
rect 355232 3742 355284 3748
rect 355244 480 355272 3742
rect 356348 480 356376 8910
rect 357544 480 357572 11834
rect 358096 3330 358124 69634
rect 359292 64874 359320 71862
rect 359464 69080 359516 69086
rect 359464 69022 359516 69028
rect 358832 64846 359320 64874
rect 358832 9110 358860 64846
rect 358820 9104 358872 9110
rect 358820 9046 358872 9052
rect 359476 8974 359504 69022
rect 360212 13122 360240 71862
rect 361592 70038 361620 71862
rect 361580 70032 361632 70038
rect 361580 69974 361632 69980
rect 362224 69760 362276 69766
rect 362224 69702 362276 69708
rect 360844 69148 360896 69154
rect 360844 69090 360896 69096
rect 360200 13116 360252 13122
rect 360200 13058 360252 13064
rect 359464 8968 359516 8974
rect 359464 8910 359516 8916
rect 359924 4820 359976 4826
rect 359924 4762 359976 4768
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 358084 3324 358136 3330
rect 358084 3266 358136 3272
rect 358740 480 358768 3606
rect 359936 480 359964 4762
rect 360856 3670 360884 69090
rect 362236 3738 362264 69702
rect 362420 69086 362448 71862
rect 362972 71862 363230 71890
rect 364030 71890 364058 72148
rect 364858 71890 364886 72148
rect 364030 71862 364104 71890
rect 362408 69080 362460 69086
rect 362408 69022 362460 69028
rect 362972 4826 363000 71862
rect 364076 69698 364104 71862
rect 364444 71862 364886 71890
rect 365686 71890 365714 72148
rect 366514 71890 366542 72148
rect 367100 71936 367152 71942
rect 365686 71862 365760 71890
rect 366514 71862 366588 71890
rect 367342 71890 367370 72148
rect 368170 71942 368198 72148
rect 367100 71878 367152 71884
rect 364064 69692 364116 69698
rect 364064 69634 364116 69640
rect 363604 69080 363656 69086
rect 363604 69022 363656 69028
rect 363616 10470 363644 69022
rect 363604 10464 363656 10470
rect 363604 10406 363656 10412
rect 364444 10402 364472 71862
rect 365732 22778 365760 71862
rect 366560 69086 366588 71862
rect 366548 69080 366600 69086
rect 366548 69022 366600 69028
rect 367112 25566 367140 71878
rect 367296 71862 367370 71890
rect 368158 71936 368210 71942
rect 368158 71878 368210 71884
rect 368998 71890 369026 72148
rect 369826 71890 369854 72148
rect 370654 71890 370682 72148
rect 371482 71890 371510 72148
rect 372310 71890 372338 72148
rect 373138 71890 373166 72148
rect 368998 71862 369072 71890
rect 369826 71862 370084 71890
rect 370654 71862 370728 71890
rect 367100 25560 367152 25566
rect 367100 25502 367152 25508
rect 365720 22772 365772 22778
rect 365720 22714 365772 22720
rect 367296 11830 367324 71862
rect 369044 69834 369072 71862
rect 369032 69828 369084 69834
rect 369032 69770 369084 69776
rect 369124 69080 369176 69086
rect 369124 69022 369176 69028
rect 367744 14476 367796 14482
rect 367744 14418 367796 14424
rect 364616 11824 364668 11830
rect 364616 11766 364668 11772
rect 367284 11824 367336 11830
rect 367284 11766 367336 11772
rect 364432 10396 364484 10402
rect 364432 10338 364484 10344
rect 363512 10328 363564 10334
rect 363512 10270 363564 10276
rect 362960 4820 363012 4826
rect 362960 4762 363012 4768
rect 361120 3732 361172 3738
rect 361120 3674 361172 3680
rect 362224 3732 362276 3738
rect 362224 3674 362276 3680
rect 360844 3664 360896 3670
rect 360844 3606 360896 3612
rect 361132 480 361160 3674
rect 362316 3528 362368 3534
rect 362316 3470 362368 3476
rect 362328 480 362356 3470
rect 363524 480 363552 10270
rect 364628 480 364656 11766
rect 367008 4956 367060 4962
rect 367008 4898 367060 4904
rect 365812 3324 365864 3330
rect 365812 3266 365864 3272
rect 365824 480 365852 3266
rect 367020 480 367048 4898
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 14418
rect 369136 3534 369164 69022
rect 370056 6322 370084 71862
rect 370700 68406 370728 71862
rect 371252 71862 371510 71890
rect 371620 71862 372338 71890
rect 372632 71862 373166 71890
rect 373966 71890 373994 72148
rect 374794 71890 374822 72148
rect 373966 71862 374040 71890
rect 370688 68400 370740 68406
rect 370688 68342 370740 68348
rect 370596 6452 370648 6458
rect 370596 6394 370648 6400
rect 370044 6316 370096 6322
rect 370044 6258 370096 6264
rect 369124 3528 369176 3534
rect 369124 3470 369176 3476
rect 369400 3460 369452 3466
rect 369400 3402 369452 3408
rect 369412 480 369440 3402
rect 370608 480 370636 6394
rect 371252 3466 371280 71862
rect 371332 13388 371384 13394
rect 371332 13330 371384 13336
rect 371240 3460 371292 3466
rect 371240 3402 371292 3408
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371344 354 371372 13330
rect 371620 13258 371648 71862
rect 372632 18698 372660 71862
rect 374012 69970 374040 71862
rect 374104 71862 374822 71890
rect 375622 71890 375650 72148
rect 376450 71890 376478 72148
rect 377278 71890 377306 72148
rect 375622 71862 375696 71890
rect 376450 71862 376524 71890
rect 374000 69964 374052 69970
rect 374000 69906 374052 69912
rect 372620 18692 372672 18698
rect 372620 18634 372672 18640
rect 374104 16574 374132 71862
rect 374644 69896 374696 69902
rect 374644 69838 374696 69844
rect 374104 16546 374224 16574
rect 371608 13252 371660 13258
rect 371608 13194 371660 13200
rect 374196 6254 374224 16546
rect 374184 6248 374236 6254
rect 374184 6190 374236 6196
rect 374092 6180 374144 6186
rect 374092 6122 374144 6128
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 374104 480 374132 6122
rect 374656 3330 374684 69838
rect 375668 66910 375696 71862
rect 376496 69902 376524 71862
rect 376864 71862 377306 71890
rect 378106 71890 378134 72148
rect 378934 71890 378962 72148
rect 379762 71890 379790 72148
rect 380590 71890 380618 72148
rect 381418 71890 381446 72148
rect 378106 71862 378180 71890
rect 376484 69896 376536 69902
rect 376484 69838 376536 69844
rect 375656 66904 375708 66910
rect 375656 66846 375708 66852
rect 376864 7614 376892 71862
rect 377404 70100 377456 70106
rect 377404 70042 377456 70048
rect 376852 7608 376904 7614
rect 376852 7550 376904 7556
rect 375288 4888 375340 4894
rect 375288 4830 375340 4836
rect 374644 3324 374696 3330
rect 374644 3266 374696 3272
rect 375300 480 375328 4830
rect 377416 3602 377444 70042
rect 378152 21418 378180 71862
rect 378244 71862 378962 71890
rect 379532 71862 379790 71890
rect 379900 71862 380618 71890
rect 380912 71862 381446 71890
rect 382246 71890 382274 72148
rect 383074 71890 383102 72148
rect 383902 72026 383930 72148
rect 383902 71998 383976 72026
rect 382246 71862 382320 71890
rect 378140 21412 378192 21418
rect 378140 21354 378192 21360
rect 378244 10334 378272 71862
rect 378416 15904 378468 15910
rect 378416 15846 378468 15852
rect 378232 10328 378284 10334
rect 378232 10270 378284 10276
rect 377680 7812 377732 7818
rect 377680 7754 377732 7760
rect 376484 3596 376536 3602
rect 376484 3538 376536 3544
rect 377404 3596 377456 3602
rect 377404 3538 377456 3544
rect 376496 480 376524 3538
rect 377692 480 377720 7754
rect 371670 354 371782 480
rect 371344 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 15846
rect 379532 7682 379560 71862
rect 379900 64874 379928 71862
rect 379624 64846 379928 64874
rect 379624 44878 379652 64846
rect 379612 44872 379664 44878
rect 379612 44814 379664 44820
rect 379520 7676 379572 7682
rect 379520 7618 379572 7624
rect 380912 3942 380940 71862
rect 382292 9042 382320 71862
rect 382384 71862 383102 71890
rect 382384 28286 382412 71862
rect 382924 70032 382976 70038
rect 382924 69974 382976 69980
rect 382372 28280 382424 28286
rect 382372 28222 382424 28228
rect 382372 11756 382424 11762
rect 382372 11698 382424 11704
rect 382280 9036 382332 9042
rect 382280 8978 382332 8984
rect 381176 7744 381228 7750
rect 381176 7686 381228 7692
rect 380900 3936 380952 3942
rect 380900 3878 380952 3884
rect 379980 3324 380032 3330
rect 379980 3266 380032 3272
rect 379992 480 380020 3266
rect 381188 480 381216 7686
rect 382384 480 382412 11698
rect 382936 3738 382964 69974
rect 383948 68338 383976 71998
rect 384730 71890 384758 72148
rect 385558 71890 385586 72148
rect 384040 71862 384758 71890
rect 385144 71862 385586 71890
rect 386386 71890 386414 72148
rect 387214 71890 387242 72148
rect 388042 71890 388070 72148
rect 388870 71890 388898 72148
rect 389698 71890 389726 72148
rect 386386 71862 386460 71890
rect 383936 68332 383988 68338
rect 383936 68274 383988 68280
rect 384040 64874 384068 71862
rect 385040 69760 385092 69766
rect 385040 69702 385092 69708
rect 383672 64846 384068 64874
rect 383672 17270 383700 64846
rect 383660 17264 383712 17270
rect 383660 17206 383712 17212
rect 384764 8968 384816 8974
rect 384764 8910 384816 8916
rect 382924 3732 382976 3738
rect 382924 3674 382976 3680
rect 383568 3664 383620 3670
rect 383568 3606 383620 3612
rect 383580 480 383608 3606
rect 384776 480 384804 8910
rect 385052 6914 385080 69702
rect 385144 8974 385172 71862
rect 385132 8968 385184 8974
rect 385132 8910 385184 8916
rect 385052 6886 386000 6914
rect 385972 480 386000 6886
rect 386432 3874 386460 71862
rect 386524 71862 387242 71890
rect 387812 71862 388070 71890
rect 388180 71862 388898 71890
rect 389192 71862 389726 71890
rect 390526 71890 390554 72148
rect 391354 71890 391382 72148
rect 392182 71890 392210 72148
rect 393010 71890 393038 72148
rect 390526 71862 390600 71890
rect 386524 14618 386552 71862
rect 386512 14612 386564 14618
rect 386512 14554 386564 14560
rect 387812 13190 387840 71862
rect 387800 13184 387852 13190
rect 387800 13126 387852 13132
rect 388180 6186 388208 71862
rect 389192 15910 389220 71862
rect 390572 31074 390600 71862
rect 390664 71862 391382 71890
rect 391952 71862 392210 71890
rect 392320 71862 393038 71890
rect 393838 71890 393866 72148
rect 394666 71890 394694 72148
rect 395494 71890 395522 72148
rect 396322 71890 396350 72148
rect 397150 71890 397178 72148
rect 393838 71862 393912 71890
rect 394666 71862 394740 71890
rect 390560 31068 390612 31074
rect 390560 31010 390612 31016
rect 389180 15904 389232 15910
rect 389180 15846 389232 15852
rect 389456 13116 389508 13122
rect 389456 13058 389508 13064
rect 388260 9104 388312 9110
rect 388260 9046 388312 9052
rect 388168 6180 388220 6186
rect 388168 6122 388220 6128
rect 386420 3868 386472 3874
rect 386420 3810 386472 3816
rect 387156 3596 387208 3602
rect 387156 3538 387208 3544
rect 387168 480 387196 3538
rect 388272 480 388300 9046
rect 389468 480 389496 13058
rect 390664 3806 390692 71862
rect 391204 69692 391256 69698
rect 391204 69634 391256 69640
rect 391112 10464 391164 10470
rect 391112 10406 391164 10412
rect 390652 3800 390704 3806
rect 390652 3742 390704 3748
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 390664 480 390692 3606
rect 391124 3482 391152 10406
rect 391216 3738 391244 69634
rect 391952 11762 391980 71862
rect 392320 64874 392348 71862
rect 393884 69698 393912 71862
rect 393964 69828 394016 69834
rect 393964 69770 394016 69776
rect 393872 69692 393924 69698
rect 393872 69634 393924 69640
rect 392044 64846 392348 64874
rect 392044 18630 392072 64846
rect 392032 18624 392084 18630
rect 392032 18566 392084 18572
rect 391940 11756 391992 11762
rect 391940 11698 391992 11704
rect 393044 4820 393096 4826
rect 393044 4762 393096 4768
rect 391204 3732 391256 3738
rect 391204 3674 391256 3680
rect 391124 3454 391888 3482
rect 391860 480 391888 3454
rect 393056 480 393084 4762
rect 393976 2990 394004 69770
rect 394712 5370 394740 71862
rect 394804 71862 395522 71890
rect 396092 71862 396350 71890
rect 396552 71862 397178 71890
rect 397978 71890 398006 72148
rect 398806 71890 398834 72148
rect 399634 71890 399662 72148
rect 400462 71890 400490 72148
rect 401290 71890 401318 72148
rect 397978 71862 398052 71890
rect 398806 71862 398880 71890
rect 394804 14482 394832 71862
rect 394792 14476 394844 14482
rect 394792 14418 394844 14424
rect 395344 10396 395396 10402
rect 395344 10338 395396 10344
rect 394700 5364 394752 5370
rect 394700 5306 394752 5312
rect 394240 3732 394292 3738
rect 394240 3674 394292 3680
rect 393964 2984 394016 2990
rect 393964 2926 394016 2932
rect 394252 480 394280 3674
rect 395356 480 395384 10338
rect 396092 3738 396120 71862
rect 396552 64874 396580 71862
rect 398024 69086 398052 71862
rect 398104 69964 398156 69970
rect 398104 69906 398156 69912
rect 398012 69080 398064 69086
rect 398012 69022 398064 69028
rect 396184 64846 396580 64874
rect 396184 5302 396212 64846
rect 396264 22772 396316 22778
rect 396264 22714 396316 22720
rect 396172 5296 396224 5302
rect 396172 5238 396224 5244
rect 396080 3732 396132 3738
rect 396080 3674 396132 3680
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396276 354 396304 22714
rect 398116 4010 398144 69906
rect 398852 69766 398880 71862
rect 398944 71862 399662 71890
rect 400232 71862 400490 71890
rect 400600 71862 401318 71890
rect 402118 71890 402146 72148
rect 402946 71890 402974 72148
rect 403774 71890 403802 72148
rect 404602 71890 404630 72148
rect 405430 71890 405458 72148
rect 406258 71890 406286 72148
rect 402118 71862 402192 71890
rect 402946 71862 403112 71890
rect 403774 71862 403848 71890
rect 398840 69760 398892 69766
rect 398840 69702 398892 69708
rect 398840 25560 398892 25566
rect 398840 25502 398892 25508
rect 398104 4004 398156 4010
rect 398104 3946 398156 3952
rect 398852 3534 398880 25502
rect 398944 5234 398972 71862
rect 399484 69080 399536 69086
rect 399484 69022 399536 69028
rect 399496 17406 399524 69022
rect 400232 46238 400260 71862
rect 400220 46232 400272 46238
rect 400220 46174 400272 46180
rect 399484 17400 399536 17406
rect 399484 17342 399536 17348
rect 399024 11824 399076 11830
rect 399024 11766 399076 11772
rect 398932 5228 398984 5234
rect 398932 5170 398984 5176
rect 397736 3528 397788 3534
rect 397736 3470 397788 3476
rect 398840 3528 398892 3534
rect 399036 3482 399064 11766
rect 400600 3670 400628 71862
rect 400864 69896 400916 69902
rect 400864 69838 400916 69844
rect 400588 3664 400640 3670
rect 400588 3606 400640 3612
rect 400876 3534 400904 69838
rect 402164 65550 402192 71862
rect 402980 68400 403032 68406
rect 402980 68342 403032 68348
rect 402152 65544 402204 65550
rect 402152 65486 402204 65492
rect 402992 6914 403020 68342
rect 403084 13122 403112 71862
rect 403820 69834 403848 71862
rect 404372 71862 404630 71890
rect 404832 71862 405458 71890
rect 405752 71862 406286 71890
rect 407086 71890 407114 72148
rect 407914 71890 407942 72148
rect 407086 71862 407160 71890
rect 403808 69828 403860 69834
rect 403808 69770 403860 69776
rect 403072 13116 403124 13122
rect 403072 13058 403124 13064
rect 402992 6886 403664 6914
rect 402520 6316 402572 6322
rect 402520 6258 402572 6264
rect 398840 3470 398892 3476
rect 397748 480 397776 3470
rect 398944 3454 399064 3482
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400864 3528 400916 3534
rect 400864 3470 400916 3476
rect 398944 480 398972 3454
rect 400140 480 400168 3470
rect 401324 2984 401376 2990
rect 401324 2926 401376 2932
rect 401336 480 401364 2926
rect 402532 480 402560 6258
rect 403636 480 403664 6886
rect 404372 5166 404400 71862
rect 404832 64874 404860 71862
rect 404464 64846 404860 64874
rect 404464 24138 404492 64846
rect 404452 24132 404504 24138
rect 404452 24074 404504 24080
rect 404360 5160 404412 5166
rect 404360 5102 404412 5108
rect 405752 3602 405780 71862
rect 406016 13252 406068 13258
rect 406016 13194 406068 13200
rect 405740 3596 405792 3602
rect 405740 3538 405792 3544
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 404832 480 404860 3402
rect 406028 480 406056 13194
rect 407132 5098 407160 71862
rect 407224 71862 407942 71890
rect 408742 71890 408770 72148
rect 409570 71890 409598 72148
rect 410398 71890 410426 72148
rect 408742 71862 408816 71890
rect 407224 25566 407252 71862
rect 408788 70038 408816 71862
rect 408880 71862 409598 71890
rect 409984 71862 410426 71890
rect 411226 71890 411254 72148
rect 412054 71890 412082 72148
rect 411226 71862 411300 71890
rect 408776 70032 408828 70038
rect 408776 69974 408828 69980
rect 407212 25560 407264 25566
rect 407212 25502 407264 25508
rect 407212 18692 407264 18698
rect 407212 18634 407264 18640
rect 407120 5092 407172 5098
rect 407120 5034 407172 5040
rect 407224 480 407252 18634
rect 408880 5030 408908 71862
rect 409880 66904 409932 66910
rect 409880 66846 409932 66852
rect 409892 16574 409920 66846
rect 409984 26926 410012 71862
rect 411272 69902 411300 71862
rect 411364 71862 412082 71890
rect 412640 71936 412692 71942
rect 412882 71890 412910 72148
rect 413710 71942 413738 72148
rect 412640 71878 412692 71884
rect 411260 69896 411312 69902
rect 411260 69838 411312 69844
rect 409972 26920 410024 26926
rect 409972 26862 410024 26868
rect 409892 16546 410840 16574
rect 409604 6248 409656 6254
rect 409604 6190 409656 6196
rect 408868 5024 408920 5030
rect 408868 4966 408920 4972
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 408420 480 408448 3946
rect 409616 480 409644 6190
rect 410812 480 410840 16546
rect 411364 4962 411392 71862
rect 411352 4956 411404 4962
rect 411352 4898 411404 4904
rect 412652 3534 412680 71878
rect 412744 71862 412910 71890
rect 413698 71936 413750 71942
rect 414538 71890 414566 72148
rect 413698 71878 413750 71884
rect 414032 71862 414566 71890
rect 415366 71890 415394 72148
rect 416194 71890 416222 72148
rect 417022 71890 417050 72148
rect 417850 71890 417878 72148
rect 418678 71890 418706 72148
rect 415366 71862 415440 71890
rect 416194 71862 416268 71890
rect 412744 29646 412772 71862
rect 412732 29640 412784 29646
rect 412732 29582 412784 29588
rect 413100 7608 413152 7614
rect 413100 7550 413152 7556
rect 411904 3528 411956 3534
rect 411904 3470 411956 3476
rect 412640 3528 412692 3534
rect 412640 3470 412692 3476
rect 411916 480 411944 3470
rect 413112 480 413140 7550
rect 414032 4894 414060 71862
rect 415412 55894 415440 71862
rect 416240 70106 416268 71862
rect 416792 71862 417050 71890
rect 417160 71862 417878 71890
rect 418264 71862 418706 71890
rect 419506 71890 419534 72148
rect 420334 71890 420362 72148
rect 421162 72026 421190 72148
rect 421162 71998 421236 72026
rect 419506 71862 419580 71890
rect 416228 70100 416280 70106
rect 416228 70042 416280 70048
rect 415400 55888 415452 55894
rect 415400 55830 415452 55836
rect 414112 21412 414164 21418
rect 414112 21354 414164 21360
rect 414124 16574 414152 21354
rect 414124 16546 414336 16574
rect 414020 4888 414072 4894
rect 414020 4830 414072 4836
rect 414308 480 414336 16546
rect 415492 10328 415544 10334
rect 415492 10270 415544 10276
rect 415504 480 415532 10270
rect 416688 7676 416740 7682
rect 416688 7618 416740 7624
rect 416700 480 416728 7618
rect 416792 4826 416820 71862
rect 416872 44872 416924 44878
rect 416872 44814 416924 44820
rect 416884 16574 416912 44814
rect 417160 32502 417188 71862
rect 417148 32496 417200 32502
rect 417148 32438 417200 32444
rect 416884 16546 417464 16574
rect 416780 4820 416832 4826
rect 416780 4762 416832 4768
rect 396510 354 396622 480
rect 396276 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418264 3466 418292 71862
rect 419552 21418 419580 71862
rect 419644 71862 420362 71890
rect 419644 42090 419672 71862
rect 421208 69970 421236 71998
rect 421990 71890 422018 72148
rect 422818 71890 422846 72148
rect 421576 71862 422018 71890
rect 422404 71862 422846 71890
rect 423646 71890 423674 72148
rect 424474 71890 424502 72148
rect 425302 71890 425330 72148
rect 426130 71890 426158 72148
rect 426958 71890 426986 72148
rect 423646 71862 423720 71890
rect 421196 69964 421248 69970
rect 421196 69906 421248 69912
rect 421576 64874 421604 71862
rect 422300 68332 422352 68338
rect 422300 68274 422352 68280
rect 420932 64846 421604 64874
rect 419632 42084 419684 42090
rect 419632 42026 419684 42032
rect 420932 22846 420960 64846
rect 421012 28280 421064 28286
rect 421012 28222 421064 28228
rect 420920 22840 420972 22846
rect 420920 22782 420972 22788
rect 419540 21412 419592 21418
rect 419540 21354 419592 21360
rect 420184 9036 420236 9042
rect 420184 8978 420236 8984
rect 418988 3936 419040 3942
rect 418988 3878 419040 3884
rect 418252 3460 418304 3466
rect 418252 3402 418304 3408
rect 419000 480 419028 3878
rect 420196 480 420224 8978
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421024 354 421052 28222
rect 422312 6914 422340 68274
rect 422404 14550 422432 71862
rect 423692 39438 423720 71862
rect 423876 71862 424502 71890
rect 425072 71862 425330 71890
rect 425440 71862 426158 71890
rect 426452 71862 426986 71890
rect 427786 71890 427814 72148
rect 428614 71890 428642 72148
rect 429442 71890 429470 72148
rect 430270 71890 430298 72148
rect 431098 71890 431126 72148
rect 427786 71862 427860 71890
rect 423680 39432 423732 39438
rect 423680 39374 423732 39380
rect 423680 17264 423732 17270
rect 423680 17206 423732 17212
rect 423692 16574 423720 17206
rect 423692 16546 423812 16574
rect 422392 14544 422444 14550
rect 422392 14486 422444 14492
rect 422312 6886 422616 6914
rect 422588 480 422616 6886
rect 423784 480 423812 16546
rect 423876 7614 423904 71862
rect 425072 28286 425100 71862
rect 425440 64874 425468 71862
rect 425164 64846 425468 64874
rect 425164 49094 425192 64846
rect 425152 49088 425204 49094
rect 425152 49030 425204 49036
rect 425060 28280 425112 28286
rect 425060 28222 425112 28228
rect 426452 9042 426480 71862
rect 427832 15978 427860 71862
rect 427924 71862 428642 71890
rect 429212 71862 429470 71890
rect 429856 71862 430298 71890
rect 430592 71862 431126 71890
rect 431926 71890 431954 72148
rect 432754 71890 432782 72148
rect 433582 71890 433610 72148
rect 431926 71862 432000 71890
rect 427924 33794 427952 71862
rect 427912 33788 427964 33794
rect 427912 33730 427964 33736
rect 427820 15972 427872 15978
rect 427820 15914 427872 15920
rect 426808 14612 426860 14618
rect 426808 14554 426860 14560
rect 426440 9036 426492 9042
rect 426440 8978 426492 8984
rect 424968 8968 425020 8974
rect 424968 8910 425020 8916
rect 423864 7608 423916 7614
rect 423864 7550 423916 7556
rect 424980 480 425008 8910
rect 426164 3868 426216 3874
rect 426164 3810 426216 3816
rect 426176 480 426204 3810
rect 421350 354 421462 480
rect 421024 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 14554
rect 428464 13184 428516 13190
rect 428464 13126 428516 13132
rect 428476 480 428504 13126
rect 429212 10402 429240 71862
rect 429856 64874 429884 71862
rect 429304 64846 429884 64874
rect 429304 57322 429332 64846
rect 429292 57316 429344 57322
rect 429292 57258 429344 57264
rect 430592 35222 430620 71862
rect 431972 44946 432000 71862
rect 432064 71862 432782 71890
rect 433352 71862 433610 71890
rect 434410 71890 434438 72148
rect 435238 71890 435266 72148
rect 434410 71862 434484 71890
rect 431960 44940 432012 44946
rect 431960 44882 432012 44888
rect 432064 38010 432092 71862
rect 433352 54602 433380 71862
rect 434456 68406 434484 71862
rect 434732 71862 435266 71890
rect 436066 71890 436094 72148
rect 436894 71890 436922 72148
rect 437722 71890 437750 72148
rect 436066 71862 436140 71890
rect 434444 68400 434496 68406
rect 434444 68342 434496 68348
rect 433340 54596 433392 54602
rect 433340 54538 433392 54544
rect 432052 38004 432104 38010
rect 432052 37946 432104 37952
rect 430580 35216 430632 35222
rect 430580 35158 430632 35164
rect 432052 31068 432104 31074
rect 432052 31010 432104 31016
rect 430856 15904 430908 15910
rect 430856 15846 430908 15852
rect 429200 10396 429252 10402
rect 429200 10338 429252 10344
rect 429660 6180 429712 6186
rect 429660 6122 429712 6128
rect 429672 480 429700 6122
rect 430868 480 430896 15846
rect 432064 480 432092 31010
rect 433984 11756 434036 11762
rect 433984 11698 434036 11704
rect 433248 3800 433300 3806
rect 433248 3742 433300 3748
rect 433260 480 433288 3742
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 11698
rect 434732 6662 434760 71862
rect 435364 69692 435416 69698
rect 435364 69634 435416 69640
rect 434812 18624 434864 18630
rect 434812 18566 434864 18572
rect 434824 16574 434852 18566
rect 434824 16546 435128 16574
rect 434720 6656 434772 6662
rect 434720 6598 434772 6604
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 435376 3398 435404 69634
rect 436112 43518 436140 71862
rect 436204 71862 436922 71890
rect 437492 71862 437750 71890
rect 438550 71890 438578 72148
rect 439378 71890 439406 72148
rect 438550 71862 438624 71890
rect 436100 43512 436152 43518
rect 436100 43454 436152 43460
rect 436204 40730 436232 71862
rect 436744 69760 436796 69766
rect 436744 69702 436796 69708
rect 436192 40724 436244 40730
rect 436192 40666 436244 40672
rect 436756 4146 436784 69702
rect 437492 6594 437520 71862
rect 438596 69086 438624 71862
rect 438964 71862 439406 71890
rect 440206 71890 440234 72148
rect 441034 71890 441062 72148
rect 440206 71862 440280 71890
rect 438584 69080 438636 69086
rect 438584 69022 438636 69028
rect 438964 11762 438992 71862
rect 439504 69080 439556 69086
rect 439504 69022 439556 69028
rect 439516 50386 439544 69022
rect 439504 50380 439556 50386
rect 439504 50322 439556 50328
rect 439136 14476 439188 14482
rect 439136 14418 439188 14424
rect 438952 11756 439004 11762
rect 438952 11698 439004 11704
rect 437480 6588 437532 6594
rect 437480 6530 437532 6536
rect 437940 5364 437992 5370
rect 437940 5306 437992 5312
rect 436744 4140 436796 4146
rect 436744 4082 436796 4088
rect 435364 3392 435416 3398
rect 435364 3334 435416 3340
rect 436744 3392 436796 3398
rect 436744 3334 436796 3340
rect 436756 480 436784 3334
rect 437952 480 437980 5306
rect 439148 480 439176 14418
rect 440252 6526 440280 71862
rect 440344 71862 441062 71890
rect 441620 71936 441672 71942
rect 441862 71890 441890 72148
rect 442690 71942 442718 72148
rect 441620 71878 441672 71884
rect 440344 51746 440372 71862
rect 440884 69828 440936 69834
rect 440884 69770 440936 69776
rect 440332 51740 440384 51746
rect 440332 51682 440384 51688
rect 440240 6520 440292 6526
rect 440240 6462 440292 6468
rect 440896 3874 440924 69770
rect 441632 6390 441660 71878
rect 441816 71862 441890 71890
rect 442678 71936 442730 71942
rect 442678 71878 442730 71884
rect 443518 71890 443546 72148
rect 444346 71890 444374 72148
rect 445174 71890 445202 72148
rect 446002 72026 446030 72148
rect 443518 71862 443592 71890
rect 444346 71862 444420 71890
rect 441712 17400 441764 17406
rect 441712 17342 441764 17348
rect 441724 16574 441752 17342
rect 441816 17270 441844 71862
rect 443564 69086 443592 71862
rect 443644 70032 443696 70038
rect 443644 69974 443696 69980
rect 443552 69080 443604 69086
rect 443552 69022 443604 69028
rect 441804 17264 441856 17270
rect 441804 17206 441856 17212
rect 441724 16546 442672 16574
rect 441620 6384 441672 6390
rect 441620 6326 441672 6332
rect 441528 5296 441580 5302
rect 441528 5238 441580 5244
rect 440884 3868 440936 3874
rect 440884 3810 440936 3816
rect 440332 3732 440384 3738
rect 440332 3674 440384 3680
rect 440344 480 440372 3674
rect 441540 480 441568 5238
rect 442644 480 442672 16546
rect 443656 3806 443684 69974
rect 444392 62898 444420 71862
rect 444484 71862 445202 71890
rect 445772 71998 446030 72026
rect 444380 62892 444432 62898
rect 444380 62834 444432 62840
rect 444484 6458 444512 71862
rect 445772 69834 445800 71998
rect 446830 71890 446858 72148
rect 447658 71890 447686 72148
rect 445864 71862 446858 71890
rect 447152 71862 447686 71890
rect 448486 71890 448514 72148
rect 449314 71890 449342 72148
rect 450142 71890 450170 72148
rect 450970 71890 450998 72148
rect 451798 71890 451826 72148
rect 448486 71862 448560 71890
rect 445760 69828 445812 69834
rect 445760 69770 445812 69776
rect 445024 69080 445076 69086
rect 445024 69022 445076 69028
rect 445036 36582 445064 69022
rect 445864 46238 445892 71862
rect 446404 69896 446456 69902
rect 446404 69838 446456 69844
rect 445760 46232 445812 46238
rect 445760 46174 445812 46180
rect 445852 46232 445904 46238
rect 445852 46174 445904 46180
rect 445024 36576 445076 36582
rect 445024 36518 445076 36524
rect 444472 6452 444524 6458
rect 444472 6394 444524 6400
rect 445024 5228 445076 5234
rect 445024 5170 445076 5176
rect 443828 4140 443880 4146
rect 443828 4082 443880 4088
rect 443644 3800 443696 3806
rect 443644 3742 443696 3748
rect 443840 480 443868 4082
rect 445036 480 445064 5170
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 46174
rect 446416 3738 446444 69838
rect 447152 6254 447180 71862
rect 448532 69698 448560 71862
rect 448624 71862 449342 71890
rect 449912 71862 450170 71890
rect 450372 71862 450998 71890
rect 451292 71862 451826 71890
rect 452626 71890 452654 72148
rect 453454 71890 453482 72148
rect 454282 71890 454310 72148
rect 455110 71890 455138 72148
rect 452626 71862 452700 71890
rect 453454 71862 453528 71890
rect 448520 69692 448572 69698
rect 448520 69634 448572 69640
rect 448520 65544 448572 65550
rect 448520 65486 448572 65492
rect 448532 6914 448560 65486
rect 448624 7682 448652 71862
rect 449808 13116 449860 13122
rect 449808 13058 449860 13064
rect 448612 7676 448664 7682
rect 448612 7618 448664 7624
rect 448532 6886 448652 6914
rect 447140 6248 447192 6254
rect 447140 6190 447192 6196
rect 446404 3732 446456 3738
rect 446404 3674 446456 3680
rect 447416 3664 447468 3670
rect 447416 3606 447468 3612
rect 447428 480 447456 3606
rect 448624 480 448652 6886
rect 449820 480 449848 13058
rect 449912 6322 449940 71862
rect 450372 64874 450400 71862
rect 450544 70100 450596 70106
rect 450544 70042 450596 70048
rect 450004 64846 450400 64874
rect 450004 49026 450032 64846
rect 449992 49020 450044 49026
rect 449992 48962 450044 48968
rect 449900 6316 449952 6322
rect 449900 6258 449952 6264
rect 450556 3670 450584 70042
rect 451292 18630 451320 71862
rect 451280 18624 451332 18630
rect 451280 18566 451332 18572
rect 452672 6186 452700 71862
rect 453500 69902 453528 71862
rect 454052 71862 454310 71890
rect 454696 71862 455138 71890
rect 455938 71890 455966 72148
rect 456766 71890 456794 72148
rect 457594 71890 457622 72148
rect 458422 72026 458450 72148
rect 458422 71998 458496 72026
rect 455938 71862 456012 71890
rect 456766 71862 456840 71890
rect 453488 69896 453540 69902
rect 453488 69838 453540 69844
rect 453304 69828 453356 69834
rect 453304 69770 453356 69776
rect 453316 32434 453344 69770
rect 453304 32428 453356 32434
rect 453304 32370 453356 32376
rect 452752 24132 452804 24138
rect 452752 24074 452804 24080
rect 452764 16574 452792 24074
rect 452764 16546 453344 16574
rect 452660 6180 452712 6186
rect 452660 6122 452712 6128
rect 452108 5160 452160 5166
rect 452108 5102 452160 5108
rect 450912 3868 450964 3874
rect 450912 3810 450964 3816
rect 450544 3664 450596 3670
rect 450544 3606 450596 3612
rect 450924 480 450952 3810
rect 452120 480 452148 5102
rect 453316 480 453344 16546
rect 454052 8974 454080 71862
rect 454696 64874 454724 71862
rect 455984 69086 456012 71862
rect 456064 69692 456116 69698
rect 456064 69634 456116 69640
rect 455972 69080 456024 69086
rect 455972 69022 456024 69028
rect 454144 64846 454724 64874
rect 454144 31074 454172 64846
rect 454132 31068 454184 31074
rect 454132 31010 454184 31016
rect 456076 22778 456104 69634
rect 456064 22772 456116 22778
rect 456064 22714 456116 22720
rect 454040 8968 454092 8974
rect 454040 8910 454092 8916
rect 456812 5302 456840 71862
rect 456996 71862 457622 71890
rect 456892 25560 456944 25566
rect 456892 25502 456944 25508
rect 456800 5296 456852 5302
rect 456800 5238 456852 5244
rect 455696 5092 455748 5098
rect 455696 5034 455748 5040
rect 454500 3596 454552 3602
rect 454500 3538 454552 3544
rect 454512 480 454540 3538
rect 455708 480 455736 5034
rect 456904 480 456932 25502
rect 456996 24138 457024 71862
rect 458468 69834 458496 71998
rect 459250 71890 459278 72148
rect 460078 71890 460106 72148
rect 458560 71862 459278 71890
rect 459572 71862 460106 71890
rect 460906 71890 460934 72148
rect 461734 71890 461762 72148
rect 462562 71890 462590 72148
rect 460906 71862 460980 71890
rect 458456 69828 458508 69834
rect 458456 69770 458508 69776
rect 458560 64874 458588 71862
rect 458824 69080 458876 69086
rect 458824 69022 458876 69028
rect 458192 64846 458588 64874
rect 456984 24132 457036 24138
rect 456984 24074 457036 24080
rect 458192 5166 458220 64846
rect 458836 44878 458864 69022
rect 458824 44872 458876 44878
rect 458824 44814 458876 44820
rect 459572 15910 459600 71862
rect 460952 69086 460980 71862
rect 461044 71862 461762 71890
rect 462332 71862 462590 71890
rect 463390 71890 463418 72148
rect 464218 71890 464246 72148
rect 463390 71862 463464 71890
rect 460940 69080 460992 69086
rect 460940 69022 460992 69028
rect 459652 26920 459704 26926
rect 459652 26862 459704 26868
rect 459664 16574 459692 26862
rect 459664 16546 459968 16574
rect 459560 15904 459612 15910
rect 459560 15846 459612 15852
rect 458180 5160 458232 5166
rect 458180 5102 458232 5108
rect 459192 5024 459244 5030
rect 459192 4966 459244 4972
rect 458088 3800 458140 3806
rect 458088 3742 458140 3748
rect 458100 480 458128 3742
rect 459204 480 459232 4966
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461044 5234 461072 71862
rect 462332 25566 462360 71862
rect 463436 69698 463464 71862
rect 463712 71862 464246 71890
rect 465046 71890 465074 72148
rect 465874 71890 465902 72148
rect 466702 71890 466730 72148
rect 467530 71890 467558 72148
rect 465046 71862 465120 71890
rect 465874 71862 465948 71890
rect 463424 69692 463476 69698
rect 463424 69634 463476 69640
rect 462320 25560 462372 25566
rect 462320 25502 462372 25508
rect 461032 5228 461084 5234
rect 461032 5170 461084 5176
rect 463712 5030 463740 71862
rect 465092 68338 465120 71862
rect 465920 70038 465948 71862
rect 466472 71862 466730 71890
rect 466840 71862 467558 71890
rect 468358 71890 468386 72148
rect 469186 71890 469214 72148
rect 470014 71890 470042 72148
rect 470842 72026 470870 72148
rect 470842 71998 470916 72026
rect 468358 71862 468432 71890
rect 469186 71862 469260 71890
rect 465908 70032 465960 70038
rect 465908 69974 465960 69980
rect 465080 68332 465132 68338
rect 465080 68274 465132 68280
rect 463792 29640 463844 29646
rect 463792 29582 463844 29588
rect 463804 16574 463832 29582
rect 463804 16546 464016 16574
rect 463700 5024 463752 5030
rect 463700 4966 463752 4972
rect 462780 4956 462832 4962
rect 462780 4898 462832 4904
rect 461584 3732 461636 3738
rect 461584 3674 461636 3680
rect 461596 480 461624 3674
rect 462792 480 462820 4898
rect 463988 480 464016 16546
rect 466472 5098 466500 71862
rect 466552 55888 466604 55894
rect 466552 55830 466604 55836
rect 466564 16574 466592 55830
rect 466840 26926 466868 71862
rect 468404 69766 468432 71862
rect 468392 69760 468444 69766
rect 468392 69702 468444 69708
rect 468484 69080 468536 69086
rect 468484 69022 468536 69028
rect 466828 26920 466880 26926
rect 466828 26862 466880 26868
rect 466564 16546 467512 16574
rect 466460 5092 466512 5098
rect 466460 5034 466512 5040
rect 466276 4888 466328 4894
rect 466276 4830 466328 4836
rect 465172 3528 465224 3534
rect 465172 3470 465224 3476
rect 465184 480 465212 3470
rect 466288 480 466316 4830
rect 467484 480 467512 16546
rect 468496 3738 468524 69022
rect 469232 4962 469260 71862
rect 469324 71862 470042 71890
rect 469324 58682 469352 71862
rect 470888 69086 470916 71998
rect 471670 71890 471698 72148
rect 472498 71890 472526 72148
rect 471256 71862 471698 71890
rect 471992 71862 472526 71890
rect 473326 71890 473354 72148
rect 474154 71890 474182 72148
rect 474982 71890 475010 72148
rect 473326 71862 473400 71890
rect 470876 69080 470928 69086
rect 470876 69022 470928 69028
rect 471256 64874 471284 71862
rect 470612 64846 471284 64874
rect 469312 58676 469364 58682
rect 469312 58618 469364 58624
rect 470612 13122 470640 64846
rect 470692 32496 470744 32502
rect 470692 32438 470744 32444
rect 470600 13116 470652 13122
rect 470600 13058 470652 13064
rect 469220 4956 469272 4962
rect 469220 4898 469272 4904
rect 469864 4820 469916 4826
rect 469864 4762 469916 4768
rect 468484 3732 468536 3738
rect 468484 3674 468536 3680
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 468680 480 468708 3606
rect 469876 480 469904 4762
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470704 354 470732 32438
rect 471992 29646 472020 71862
rect 472624 69080 472676 69086
rect 472624 69022 472676 69028
rect 471980 29640 472032 29646
rect 471980 29582 472032 29588
rect 472636 3670 472664 69022
rect 473372 57254 473400 71862
rect 473464 71862 474182 71890
rect 474844 71862 475010 71890
rect 475810 71890 475838 72148
rect 476638 71890 476666 72148
rect 475810 71862 475884 71890
rect 473360 57248 473412 57254
rect 473360 57190 473412 57196
rect 473360 42084 473412 42090
rect 473360 42026 473412 42032
rect 472624 3664 472676 3670
rect 472624 3606 472676 3612
rect 473372 3534 473400 42026
rect 473464 10334 473492 71862
rect 474740 69964 474792 69970
rect 474740 69906 474792 69912
rect 473544 21412 473596 21418
rect 473544 21354 473596 21360
rect 473452 10328 473504 10334
rect 473452 10270 473504 10276
rect 473556 6914 473584 21354
rect 474752 16574 474780 69906
rect 474844 21418 474872 71862
rect 475856 69086 475884 71862
rect 476132 71862 476666 71890
rect 477466 71890 477494 72148
rect 478294 71890 478322 72148
rect 479122 72026 479150 72148
rect 479122 71998 479196 72026
rect 477466 71862 477540 71890
rect 478294 71862 478368 71890
rect 475844 69080 475896 69086
rect 475844 69022 475896 69028
rect 474832 21412 474884 21418
rect 474832 21354 474884 21360
rect 474752 16546 475792 16574
rect 473464 6886 473584 6914
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 472256 3460 472308 3466
rect 472256 3402 472308 3408
rect 472268 480 472296 3402
rect 473464 480 473492 6886
rect 474188 3528 474240 3534
rect 474188 3470 474240 3476
rect 471030 354 471142 480
rect 470704 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3470
rect 475764 480 475792 16546
rect 476132 14482 476160 71862
rect 476764 69080 476816 69086
rect 476764 69022 476816 69028
rect 476776 43450 476804 69022
rect 476764 43444 476816 43450
rect 476764 43386 476816 43392
rect 477512 39370 477540 71862
rect 478144 70032 478196 70038
rect 478144 69974 478196 69980
rect 477500 39364 477552 39370
rect 477500 39306 477552 39312
rect 476212 22840 476264 22846
rect 476212 22782 476264 22788
rect 476224 16574 476252 22782
rect 478156 16574 478184 69974
rect 478340 69970 478368 71862
rect 478328 69964 478380 69970
rect 478328 69906 478380 69912
rect 479168 66910 479196 71998
rect 479950 71890 479978 72148
rect 479536 71862 479978 71890
rect 480778 71890 480806 72148
rect 481606 71890 481634 72148
rect 482434 71890 482462 72148
rect 480778 71862 480852 71890
rect 481606 71862 481680 71890
rect 479156 66904 479208 66910
rect 479156 66846 479208 66852
rect 479536 64874 479564 71862
rect 480824 69086 480852 71862
rect 480812 69080 480864 69086
rect 480812 69022 480864 69028
rect 478892 64846 479564 64874
rect 478892 62830 478920 64846
rect 481652 64190 481680 71862
rect 481744 71862 482462 71890
rect 483262 71890 483290 72148
rect 484090 71890 484118 72148
rect 484918 71890 484946 72148
rect 483262 71862 483336 71890
rect 484090 71862 484164 71890
rect 481640 64184 481692 64190
rect 481640 64126 481692 64132
rect 478880 62824 478932 62830
rect 478880 62766 478932 62772
rect 481640 49088 481692 49094
rect 481640 49030 481692 49036
rect 478880 39432 478932 39438
rect 478880 39374 478932 39380
rect 476224 16546 476528 16574
rect 478156 16546 478276 16574
rect 476120 14476 476172 14482
rect 476120 14418 476172 14424
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478144 14544 478196 14550
rect 478144 14486 478196 14492
rect 478156 480 478184 14486
rect 478248 3806 478276 16546
rect 478236 3800 478288 3806
rect 478236 3742 478288 3748
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 39374
rect 480536 7608 480588 7614
rect 480536 7550 480588 7556
rect 480548 480 480576 7550
rect 481652 3534 481680 49030
rect 481744 42090 481772 71862
rect 483308 70174 483336 71862
rect 483296 70168 483348 70174
rect 483296 70110 483348 70116
rect 482284 69080 482336 69086
rect 482284 69022 482336 69028
rect 481732 42084 481784 42090
rect 481732 42026 481784 42032
rect 481732 28280 481784 28286
rect 481732 28222 481784 28228
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 28222
rect 482296 3602 482324 69022
rect 484136 65550 484164 71862
rect 484412 71862 484946 71890
rect 485746 71890 485774 72148
rect 486574 71890 486602 72148
rect 487402 71890 487430 72148
rect 485746 71862 485820 71890
rect 484124 65544 484176 65550
rect 484124 65486 484176 65492
rect 484412 61402 484440 71862
rect 484400 61396 484452 61402
rect 484400 61338 484452 61344
rect 485792 37942 485820 71862
rect 485884 71862 486602 71890
rect 487172 71862 487430 71890
rect 488230 71890 488258 72148
rect 489058 71890 489086 72148
rect 488230 71862 488304 71890
rect 485780 37936 485832 37942
rect 485780 37878 485832 37884
rect 485780 33788 485832 33794
rect 485780 33730 485832 33736
rect 484768 15972 484820 15978
rect 484768 15914 484820 15920
rect 484032 9036 484084 9042
rect 484032 8978 484084 8984
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 8978
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 15914
rect 485792 6914 485820 33730
rect 485884 7614 485912 71862
rect 487172 55894 487200 71862
rect 488276 70106 488304 71862
rect 488552 71862 489086 71890
rect 489886 71890 489914 72148
rect 490714 71890 490742 72148
rect 491542 71890 491570 72148
rect 492370 71890 492398 72148
rect 489886 71862 489960 71890
rect 488264 70100 488316 70106
rect 488264 70042 488316 70048
rect 487160 55888 487212 55894
rect 487160 55830 487212 55836
rect 487160 10396 487212 10402
rect 487160 10338 487212 10344
rect 485872 7608 485924 7614
rect 485872 7550 485924 7556
rect 485792 6886 486464 6914
rect 486436 480 486464 6886
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 10338
rect 488552 4826 488580 71862
rect 489932 67658 489960 71862
rect 490024 71862 490742 71890
rect 491312 71862 491570 71890
rect 491680 71862 492398 71890
rect 493198 71890 493226 72148
rect 494026 71890 494054 72148
rect 494854 71890 494882 72148
rect 495682 71890 495710 72148
rect 493198 71862 493272 71890
rect 494026 71862 494100 71890
rect 494854 71862 494928 71890
rect 489920 67652 489972 67658
rect 489920 67594 489972 67600
rect 488632 57316 488684 57322
rect 488632 57258 488684 57264
rect 488644 16574 488672 57258
rect 490024 54534 490052 71862
rect 490196 67652 490248 67658
rect 490196 67594 490248 67600
rect 490012 54528 490064 54534
rect 490012 54470 490064 54476
rect 489920 44940 489972 44946
rect 489920 44882 489972 44888
rect 488644 16546 488856 16574
rect 488540 4820 488592 4826
rect 488540 4762 488592 4768
rect 488828 480 488856 16546
rect 489932 3534 489960 44882
rect 490012 35216 490064 35222
rect 490012 35158 490064 35164
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 35158
rect 490208 33794 490236 67594
rect 490196 33788 490248 33794
rect 490196 33730 490248 33736
rect 491312 4894 491340 71862
rect 491680 64874 491708 71862
rect 493244 70174 493272 71862
rect 493232 70168 493284 70174
rect 493232 70110 493284 70116
rect 491404 64846 491708 64874
rect 491404 53106 491432 64846
rect 492680 54596 492732 54602
rect 492680 54538 492732 54544
rect 491392 53100 491444 53106
rect 491392 53042 491444 53048
rect 491392 38004 491444 38010
rect 491392 37946 491444 37952
rect 491404 16574 491432 37946
rect 492692 16574 492720 54538
rect 491404 16546 492352 16574
rect 492692 16546 493088 16574
rect 491300 4888 491352 4894
rect 491300 4830 491352 4836
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494072 3534 494100 71862
rect 494900 70242 494928 71862
rect 495544 71862 495710 71890
rect 494704 70236 494756 70242
rect 494704 70178 494756 70184
rect 494888 70236 494940 70242
rect 494888 70178 494940 70184
rect 494716 70038 494744 70178
rect 494704 70032 494756 70038
rect 494704 69974 494756 69980
rect 494152 68400 494204 68406
rect 494152 68342 494204 68348
rect 494164 16574 494192 68342
rect 494164 16546 494744 16574
rect 494060 3528 494112 3534
rect 494060 3470 494112 3476
rect 494716 480 494744 16546
rect 495544 3466 495572 71862
rect 507860 62892 507912 62898
rect 507860 62834 507912 62840
rect 503720 51740 503772 51746
rect 503720 51682 503772 51688
rect 499580 50380 499632 50386
rect 499580 50322 499632 50328
rect 496820 43512 496872 43518
rect 496820 43454 496872 43460
rect 496832 16574 496860 43454
rect 498200 40724 498252 40730
rect 498200 40666 498252 40672
rect 496832 16546 497136 16574
rect 495900 6656 495952 6662
rect 495900 6598 495952 6604
rect 495532 3460 495584 3466
rect 495532 3402 495584 3408
rect 495912 480 495940 6598
rect 497108 480 497136 16546
rect 498212 480 498240 40666
rect 499592 16574 499620 50322
rect 499592 16546 500632 16574
rect 499396 6588 499448 6594
rect 499396 6530 499448 6536
rect 499408 480 499436 6530
rect 500604 480 500632 16546
rect 501328 11756 501380 11762
rect 501328 11698 501380 11704
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 354 501368 11698
rect 502984 6520 503036 6526
rect 502984 6462 503036 6468
rect 502996 480 503024 6462
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 51682
rect 506480 36576 506532 36582
rect 506480 36518 506532 36524
rect 505100 17264 505152 17270
rect 505100 17206 505152 17212
rect 505112 16574 505140 17206
rect 506492 16574 506520 36518
rect 507872 16574 507900 62834
rect 510620 32428 510672 32434
rect 510620 32370 510672 32376
rect 510632 16574 510660 32370
rect 505112 16546 505416 16574
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511028 16574
rect 505388 480 505416 16546
rect 506480 6384 506532 6390
rect 506480 6326 506532 6332
rect 506492 480 506520 6326
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 510068 6452 510120 6458
rect 510068 6394 510120 6400
rect 510080 480 510108 6394
rect 511000 3482 511028 16546
rect 511092 6866 511120 633490
rect 511448 632868 511500 632874
rect 511448 632810 511500 632816
rect 511356 632460 511408 632466
rect 511356 632402 511408 632408
rect 511262 630728 511318 630737
rect 511262 630663 511318 630672
rect 511276 86970 511304 630663
rect 511368 206990 511396 632402
rect 511460 299470 511488 632810
rect 511448 299464 511500 299470
rect 511448 299406 511500 299412
rect 511356 206984 511408 206990
rect 511356 206926 511408 206932
rect 511264 86964 511316 86970
rect 511264 86906 511316 86912
rect 512012 20670 512040 633558
rect 512092 633480 512144 633486
rect 512092 633422 512144 633428
rect 512104 59362 512132 633422
rect 512092 59356 512144 59362
rect 512092 59298 512144 59304
rect 512656 46918 512684 634879
rect 512748 564398 512776 635326
rect 512840 618254 512868 635394
rect 512828 618248 512880 618254
rect 512828 618190 512880 618196
rect 512736 564392 512788 564398
rect 512736 564334 512788 564340
rect 512644 46912 512696 46918
rect 512644 46854 512696 46860
rect 512092 46232 512144 46238
rect 512092 46174 512144 46180
rect 512000 20664 512052 20670
rect 512000 20606 512052 20612
rect 511080 6860 511132 6866
rect 511080 6802 511132 6808
rect 511000 3454 511304 3482
rect 511276 480 511304 3454
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512104 354 512132 46174
rect 514036 33114 514064 636239
rect 514116 634840 514168 634846
rect 514116 634782 514168 634788
rect 514128 126954 514156 634782
rect 514220 167006 514248 636618
rect 514300 635248 514352 635254
rect 514300 635190 514352 635196
rect 514312 511970 514340 635190
rect 514300 511964 514352 511970
rect 514300 511906 514352 511912
rect 514208 167000 514260 167006
rect 514208 166942 514260 166948
rect 514116 126948 514168 126954
rect 514116 126890 514168 126896
rect 515416 100706 515444 637638
rect 516784 637628 516836 637634
rect 516784 637570 516836 637576
rect 516796 113150 516824 637570
rect 516968 636948 517020 636954
rect 516968 636890 517020 636896
rect 516876 636812 516928 636818
rect 516876 636754 516928 636760
rect 516888 245614 516916 636754
rect 516980 405686 517008 636890
rect 518164 633956 518216 633962
rect 518164 633898 518216 633904
rect 516968 405680 517020 405686
rect 516968 405622 517020 405628
rect 516876 245608 516928 245614
rect 516876 245550 516928 245556
rect 518176 179382 518204 633898
rect 518268 273222 518296 637842
rect 520936 325650 520964 637978
rect 521028 379506 521056 638046
rect 522304 634024 522356 634030
rect 522304 633966 522356 633972
rect 521016 379500 521068 379506
rect 521016 379442 521068 379448
rect 520924 325644 520976 325650
rect 520924 325586 520976 325592
rect 518256 273216 518308 273222
rect 518256 273158 518308 273164
rect 522316 259418 522344 633966
rect 522408 431934 522436 638182
rect 549916 637022 549944 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 549904 637016 549956 637022
rect 549904 636958 549956 636964
rect 531964 636268 532016 636274
rect 531964 636210 532016 636216
rect 525248 635112 525300 635118
rect 525248 635054 525300 635060
rect 525156 634228 525208 634234
rect 525156 634170 525208 634176
rect 525064 634092 525116 634098
rect 525064 634034 525116 634040
rect 522396 431928 522448 431934
rect 522396 431870 522448 431876
rect 525076 313274 525104 634034
rect 525168 365702 525196 634170
rect 525260 471986 525288 635054
rect 525248 471980 525300 471986
rect 525248 471922 525300 471928
rect 525156 365696 525208 365702
rect 525156 365638 525208 365644
rect 525064 313268 525116 313274
rect 525064 313210 525116 313216
rect 522304 259412 522356 259418
rect 522304 259354 522356 259360
rect 518164 179376 518216 179382
rect 518164 179318 518216 179324
rect 516784 113144 516836 113150
rect 516784 113086 516836 113092
rect 515404 100700 515456 100706
rect 515404 100642 515456 100648
rect 531976 73166 532004 636210
rect 545764 634160 545816 634166
rect 545764 634102 545816 634108
rect 545776 458182 545804 634102
rect 577870 633856 577926 633865
rect 577870 633791 577926 633800
rect 577686 633584 577742 633593
rect 577686 633519 577742 633528
rect 577502 633448 577558 633457
rect 577502 633383 577558 633392
rect 545764 458176 545816 458182
rect 545764 458118 545816 458124
rect 531964 73160 532016 73166
rect 531964 73102 532016 73108
rect 549904 70236 549956 70242
rect 549904 70178 549956 70184
rect 548524 70168 548576 70174
rect 548524 70110 548576 70116
rect 547144 70100 547196 70106
rect 547144 70042 547196 70048
rect 545764 70032 545816 70038
rect 545764 69974 545816 69980
rect 543004 69964 543056 69970
rect 543004 69906 543056 69912
rect 521660 69896 521712 69902
rect 521660 69838 521712 69844
rect 517520 49020 517572 49026
rect 517520 48962 517572 48968
rect 514024 33108 514076 33114
rect 514024 33050 514076 33056
rect 514760 22772 514812 22778
rect 514760 22714 514812 22720
rect 513564 6248 513616 6254
rect 513564 6190 513616 6196
rect 513576 480 513604 6190
rect 514772 480 514800 22714
rect 517532 16574 517560 48962
rect 518900 18624 518952 18630
rect 518900 18566 518952 18572
rect 518912 16574 518940 18566
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515956 7676 516008 7682
rect 515956 7618 516008 7624
rect 515968 480 515996 7618
rect 517152 6316 517204 6322
rect 517152 6258 517204 6264
rect 517164 480 517192 6258
rect 512430 354 512542 480
rect 512104 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 520740 6180 520792 6186
rect 520740 6122 520792 6128
rect 520752 480 520780 6122
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521672 354 521700 69838
rect 528560 69828 528612 69834
rect 528560 69770 528612 69776
rect 524420 44872 524472 44878
rect 524420 44814 524472 44820
rect 523040 31068 523092 31074
rect 523040 31010 523092 31016
rect 523052 16574 523080 31010
rect 524432 16574 524460 44814
rect 527180 24132 527232 24138
rect 527180 24074 527232 24080
rect 527192 16574 527220 24074
rect 523052 16546 523816 16574
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 523040 8968 523092 8974
rect 523040 8910 523092 8916
rect 523052 480 523080 8910
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 526628 5296 526680 5302
rect 526628 5238 526680 5244
rect 526640 480 526668 5238
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 69770
rect 540244 69760 540296 69766
rect 540244 69702 540296 69708
rect 535460 69692 535512 69698
rect 535460 69634 535512 69640
rect 534080 25560 534132 25566
rect 534080 25502 534132 25508
rect 534092 16574 534120 25502
rect 535472 16574 535500 69634
rect 538220 68332 538272 68338
rect 538220 68274 538272 68280
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 531320 15904 531372 15910
rect 531320 15846 531372 15852
rect 530124 5160 530176 5166
rect 530124 5102 530176 5108
rect 530136 480 530164 5102
rect 531332 480 531360 15846
rect 533712 5228 533764 5234
rect 533712 5170 533764 5176
rect 532516 3732 532568 3738
rect 532516 3674 532568 3680
rect 532528 480 532556 3674
rect 533724 480 533752 5170
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537208 5024 537260 5030
rect 537208 4966 537260 4972
rect 537220 480 537248 4966
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 68274
rect 539600 3800 539652 3806
rect 539600 3742 539652 3748
rect 539612 480 539640 3742
rect 540256 3194 540284 69702
rect 540980 26920 541032 26926
rect 540980 26862 541032 26868
rect 540992 16574 541020 26862
rect 540992 16546 542032 16574
rect 540796 5092 540848 5098
rect 540796 5034 540848 5040
rect 540244 3188 540296 3194
rect 540244 3130 540296 3136
rect 540808 480 540836 5034
rect 542004 480 542032 16546
rect 543016 3942 543044 69906
rect 545120 58676 545172 58682
rect 545120 58618 545172 58624
rect 545132 16574 545160 58618
rect 545132 16546 545528 16574
rect 544384 4956 544436 4962
rect 544384 4898 544436 4904
rect 543004 3936 543056 3942
rect 543004 3878 543056 3884
rect 543188 3188 543240 3194
rect 543188 3130 543240 3136
rect 543200 480 543228 3130
rect 544396 480 544424 4898
rect 545500 480 545528 16546
rect 545776 3874 545804 69974
rect 545764 3868 545816 3874
rect 545764 3810 545816 3816
rect 547156 3806 547184 70042
rect 547880 29640 547932 29646
rect 547880 29582 547932 29588
rect 547144 3800 547196 3806
rect 547144 3742 547196 3748
rect 546684 3664 546736 3670
rect 546684 3606 546736 3612
rect 546696 480 546724 3606
rect 547892 3398 547920 29582
rect 547972 13116 548024 13122
rect 547972 13058 548024 13064
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 3210 548012 13058
rect 548536 3738 548564 70110
rect 549260 57248 549312 57254
rect 549260 57190 549312 57196
rect 549272 16574 549300 57190
rect 549272 16546 549852 16574
rect 548524 3732 548576 3738
rect 548524 3674 548576 3680
rect 549824 3482 549852 16546
rect 549916 3670 549944 70178
rect 557540 66904 557592 66910
rect 557540 66846 557592 66852
rect 553400 43444 553452 43450
rect 553400 43386 553452 43392
rect 552020 21412 552072 21418
rect 552020 21354 552072 21360
rect 552032 16574 552060 21354
rect 553412 16574 553440 43386
rect 556252 39364 556304 39370
rect 556252 39306 556304 39312
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 551008 10328 551060 10334
rect 551008 10270 551060 10276
rect 549904 3664 549956 3670
rect 549904 3606 549956 3612
rect 549824 3454 550312 3482
rect 548708 3392 548760 3398
rect 548708 3334 548760 3340
rect 547892 3182 548012 3210
rect 547892 480 547920 3182
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548720 354 548748 3334
rect 550284 480 550312 3454
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 10270
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554780 14476 554832 14482
rect 554780 14418 554832 14424
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 14418
rect 556264 6914 556292 39306
rect 557552 16574 557580 66846
rect 564532 65544 564584 65550
rect 564532 65486 564584 65492
rect 561680 64184 561732 64190
rect 561680 64126 561732 64132
rect 558920 62824 558972 62830
rect 558920 62766 558972 62772
rect 558932 16574 558960 62766
rect 561692 16574 561720 64126
rect 563060 42084 563112 42090
rect 563060 42026 563112 42032
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 561692 16546 562088 16574
rect 556172 6886 556292 6914
rect 556172 480 556200 6886
rect 557356 3936 557408 3942
rect 557356 3878 557408 3884
rect 557368 480 557396 3878
rect 558564 480 558592 16546
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560852 3596 560904 3602
rect 560852 3538 560904 3544
rect 560864 480 560892 3538
rect 562060 480 562088 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 559718 -960 559830 326
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 42026
rect 564544 16574 564572 65486
rect 565820 61396 565872 61402
rect 565820 61338 565872 61344
rect 565832 16574 565860 61338
rect 569960 55888 570012 55894
rect 569960 55830 570012 55836
rect 567200 37936 567252 37942
rect 567200 37878 567252 37884
rect 567212 16574 567240 37878
rect 569972 16574 570000 55830
rect 574100 54528 574152 54534
rect 574100 54470 574152 54476
rect 572720 33788 572772 33794
rect 572720 33730 572772 33736
rect 572732 16574 572760 33730
rect 574112 16574 574140 54470
rect 576124 53100 576176 53106
rect 576124 53042 576176 53048
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 7608 569184 7614
rect 569132 7550 569184 7556
rect 569144 480 569172 7550
rect 570340 480 570368 16546
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 571524 3800 571576 3806
rect 571524 3742 571576 3748
rect 571536 480 571564 3742
rect 572732 480 572760 4762
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576136 3262 576164 53042
rect 577516 6798 577544 633383
rect 577700 20670 577728 633519
rect 577884 60722 577912 633791
rect 579988 632800 580040 632806
rect 579988 632742 580040 632748
rect 580000 630766 580028 632742
rect 580448 632732 580500 632738
rect 580448 632674 580500 632680
rect 580080 632664 580132 632670
rect 580080 632606 580132 632612
rect 579988 630760 580040 630766
rect 579988 630702 580040 630708
rect 579988 618248 580040 618254
rect 579988 618190 580040 618196
rect 580000 617545 580028 618190
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 580092 591025 580120 632606
rect 580264 632120 580316 632126
rect 580264 632062 580316 632068
rect 580172 631100 580224 631106
rect 580172 631042 580224 631048
rect 580184 630873 580212 631042
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 630760 580224 630766
rect 580172 630702 580224 630708
rect 580078 591016 580134 591025
rect 580078 590951 580134 590960
rect 580184 577697 580212 630702
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 579804 471980 579856 471986
rect 579804 471922 579856 471928
rect 579816 471481 579844 471922
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 579620 379500 579672 379506
rect 579620 379442 579672 379448
rect 579632 378457 579660 379442
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 579712 313268 579764 313274
rect 579712 313210 579764 313216
rect 579724 312089 579752 313210
rect 579710 312080 579766 312089
rect 579710 312015 579766 312024
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 298761 579844 299406
rect 579802 298752 579858 298761
rect 579802 298687 579858 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580276 192545 580304 632062
rect 580356 630692 580408 630698
rect 580356 630634 580408 630640
rect 580368 219065 580396 630634
rect 580460 232393 580488 632674
rect 580908 632528 580960 632534
rect 580908 632470 580960 632476
rect 580724 632324 580776 632330
rect 580724 632266 580776 632272
rect 580632 630964 580684 630970
rect 580632 630906 580684 630912
rect 580540 630896 580592 630902
rect 580540 630838 580592 630844
rect 580552 351937 580580 630838
rect 580644 418305 580672 630906
rect 580736 484673 580764 632266
rect 580816 631032 580868 631038
rect 580816 630974 580868 630980
rect 580828 524521 580856 630974
rect 580920 537849 580948 632470
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580630 418296 580686 418305
rect 580630 418231 580686 418240
rect 580538 351928 580594 351937
rect 580538 351863 580594 351872
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 580262 192536 580318 192545
rect 580262 192471 580318 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 577872 60716 577924 60722
rect 577872 60658 577924 60664
rect 579988 60716 580040 60722
rect 579988 60658 580040 60664
rect 580000 59673 580028 60658
rect 579986 59664 580042 59673
rect 579986 59599 580042 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 577688 20664 577740 20670
rect 577688 20606 577740 20612
rect 579804 20664 579856 20670
rect 579804 20606 579856 20612
rect 579816 19825 579844 20606
rect 579802 19816 579858 19825
rect 579802 19751 579858 19760
rect 577504 6792 577556 6798
rect 577504 6734 577556 6740
rect 579712 6792 579764 6798
rect 579712 6734 579764 6740
rect 579724 6633 579752 6734
rect 579710 6624 579766 6633
rect 579710 6559 579766 6568
rect 576308 4888 576360 4894
rect 576308 4830 576360 4836
rect 576124 3256 576176 3262
rect 576124 3198 576176 3204
rect 576320 480 576348 4830
rect 578608 3732 578660 3738
rect 578608 3674 578660 3680
rect 577412 3256 577464 3262
rect 577412 3198 577464 3204
rect 577424 480 577452 3198
rect 578620 480 578648 3674
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 582208 480 582236 3606
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3146 619112 3202 619168
rect 2778 606056 2834 606112
rect 3146 579944 3202 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 3330 527856 3386 527912
rect 3330 501780 3332 501800
rect 3332 501780 3384 501800
rect 3384 501780 3386 501800
rect 3330 501744 3386 501780
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 397432 3386 397488
rect 2778 371320 2834 371376
rect 2962 345344 3018 345400
rect 2778 319232 2834 319288
rect 3238 267144 3294 267200
rect 2778 254088 2834 254144
rect 3330 214920 3386 214976
rect 3514 632032 3570 632088
rect 3514 631216 3570 631272
rect 4066 514800 4122 514856
rect 3974 449520 4030 449576
rect 3882 358400 3938 358456
rect 3790 306176 3846 306232
rect 3698 293120 3754 293176
rect 3606 241032 3662 241088
rect 3514 201864 3570 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 2778 149776 2834 149832
rect 3422 110608 3478 110664
rect 2778 97552 2834 97608
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 82726 636248 82782 636304
rect 79138 633392 79194 633448
rect 90454 634888 90510 634944
rect 86682 633528 86738 633584
rect 97906 633800 97962 633856
rect 120630 632304 120686 632360
rect 116858 632032 116914 632088
rect 101770 631352 101826 631408
rect 467332 632168 467388 632224
rect 478326 633936 478382 633992
rect 490010 633664 490066 633720
rect 514022 636248 514078 636304
rect 512642 634888 512698 634944
rect 415490 631488 415546 631544
rect 416594 631488 416650 631544
rect 366546 631352 366602 631408
rect 410522 631388 410524 631408
rect 410524 631388 410576 631408
rect 410576 631388 410578 631408
rect 410522 631352 410578 631388
rect 417974 631352 418030 631408
rect 511262 630672 511318 630728
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 577870 633800 577926 633856
rect 577686 633528 577742 633584
rect 577502 633392 577558 633448
rect 579986 617480 580042 617536
rect 580170 630808 580226 630864
rect 580078 590960 580134 591016
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 511264 580226 511320
rect 579802 471416 579858 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 579618 378392 579674 378448
rect 580170 365064 580226 365120
rect 580170 325216 580226 325272
rect 579710 312024 579766 312080
rect 579802 298696 579858 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 205672 580226 205728
rect 580906 537784 580962 537840
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 580630 418240 580686 418296
rect 580538 351872 580594 351928
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 580262 192480 580318 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 579986 59608 580042 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579802 19760 579858 19816
rect 579710 6568 579766 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 82721 636306 82787 636309
rect 514017 636306 514083 636309
rect 82721 636304 514083 636306
rect 82721 636248 82726 636304
rect 82782 636248 514022 636304
rect 514078 636248 514083 636304
rect 82721 636246 514083 636248
rect 82721 636243 82787 636246
rect 514017 636243 514083 636246
rect 90449 634946 90515 634949
rect 512637 634946 512703 634949
rect 90449 634944 512703 634946
rect 90449 634888 90454 634944
rect 90510 634888 512642 634944
rect 512698 634888 512703 634944
rect 90449 634886 512703 634888
rect 90449 634883 90515 634886
rect 512637 634883 512703 634886
rect 3550 633932 3556 633996
rect 3620 633994 3626 633996
rect 478321 633994 478387 633997
rect 3620 633992 478387 633994
rect 3620 633936 478326 633992
rect 478382 633936 478387 633992
rect 3620 633934 478387 633936
rect 3620 633932 3626 633934
rect 478321 633931 478387 633934
rect 97901 633858 97967 633861
rect 577865 633858 577931 633861
rect 97901 633856 577931 633858
rect 97901 633800 97906 633856
rect 97962 633800 577870 633856
rect 577926 633800 577931 633856
rect 97901 633798 577931 633800
rect 97901 633795 97967 633798
rect 577865 633795 577931 633798
rect 3366 633660 3372 633724
rect 3436 633722 3442 633724
rect 490005 633722 490071 633725
rect 3436 633720 490071 633722
rect 3436 633664 490010 633720
rect 490066 633664 490071 633720
rect 3436 633662 490071 633664
rect 3436 633660 3442 633662
rect 490005 633659 490071 633662
rect 86677 633586 86743 633589
rect 577681 633586 577747 633589
rect 86677 633584 577747 633586
rect 86677 633528 86682 633584
rect 86738 633528 577686 633584
rect 577742 633528 577747 633584
rect 86677 633526 577747 633528
rect 86677 633523 86743 633526
rect 577681 633523 577747 633526
rect 79133 633450 79199 633453
rect 577497 633450 577563 633453
rect 79133 633448 140790 633450
rect 79133 633392 79138 633448
rect 79194 633392 140790 633448
rect 79133 633390 140790 633392
rect 79133 633387 79199 633390
rect 140730 633314 140790 633390
rect 150390 633390 411270 633450
rect 150390 633314 150450 633390
rect 140730 633254 150450 633314
rect 411210 633314 411270 633390
rect 420870 633448 577563 633450
rect 420870 633392 577502 633448
rect 577558 633392 577563 633448
rect 420870 633390 577563 633392
rect 420870 633314 420930 633390
rect 577497 633387 577563 633390
rect 411210 633254 420930 633314
rect 120625 632362 120691 632365
rect 580206 632362 580212 632364
rect 120625 632360 580212 632362
rect 120625 632304 120630 632360
rect 120686 632304 580212 632360
rect 120625 632302 580212 632304
rect 120625 632299 120691 632302
rect 580206 632300 580212 632302
rect 580276 632300 580282 632364
rect -960 632090 480 632180
rect 3734 632164 3740 632228
rect 3804 632226 3810 632228
rect 467327 632226 467393 632229
rect 3804 632224 467393 632226
rect 3804 632168 467332 632224
rect 467388 632168 467393 632224
rect 3804 632166 467393 632168
rect 3804 632164 3810 632166
rect 467327 632163 467393 632166
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 116853 632090 116919 632093
rect 580390 632090 580396 632092
rect 116853 632088 580396 632090
rect 116853 632032 116858 632088
rect 116914 632032 580396 632088
rect 116853 632030 580396 632032
rect 116853 632027 116919 632030
rect 580390 632028 580396 632030
rect 580460 632028 580466 632092
rect 415485 631546 415551 631549
rect 416589 631546 416655 631549
rect 415485 631544 416655 631546
rect 415485 631488 415490 631544
rect 415546 631488 416594 631544
rect 416650 631488 416655 631544
rect 415485 631486 416655 631488
rect 415485 631483 415551 631486
rect 416589 631483 416655 631486
rect 101765 631410 101831 631413
rect 108246 631410 108252 631412
rect 101765 631408 108252 631410
rect 101765 631352 101770 631408
rect 101826 631352 108252 631408
rect 101765 631350 108252 631352
rect 101765 631347 101831 631350
rect 108246 631348 108252 631350
rect 108316 631348 108322 631412
rect 366541 631410 366607 631413
rect 354630 631408 366607 631410
rect 354630 631352 366546 631408
rect 366602 631352 366607 631408
rect 354630 631350 366607 631352
rect 3509 631274 3575 631277
rect 354630 631274 354690 631350
rect 366541 631347 366607 631350
rect 410517 631410 410583 631413
rect 417969 631410 418035 631413
rect 410517 631408 418035 631410
rect 410517 631352 410522 631408
rect 410578 631352 417974 631408
rect 418030 631352 418035 631408
rect 410517 631350 418035 631352
rect 410517 631347 410583 631350
rect 417969 631347 418035 631350
rect 3509 631272 354690 631274
rect 3509 631216 3514 631272
rect 3570 631216 354690 631272
rect 3509 631214 354690 631216
rect 3509 631211 3575 631214
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 108246 630668 108252 630732
rect 108316 630730 108322 630732
rect 511257 630730 511323 630733
rect 108316 630728 511323 630730
rect 108316 630672 511262 630728
rect 511318 630672 511323 630728
rect 583520 630716 584960 630806
rect 108316 630670 511323 630672
rect 108316 630668 108322 630670
rect 511257 630667 511323 630670
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580073 591018 580139 591021
rect 583520 591018 584960 591108
rect 580073 591016 584960 591018
rect 580073 590960 580078 591016
rect 580134 590960 584960 591016
rect 580073 590958 584960 590960
rect 580073 590955 580139 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3969 449578 4035 449581
rect -960 449576 4035 449578
rect -960 449520 3974 449576
rect 4030 449520 4035 449576
rect -960 449518 4035 449520
rect -960 449428 480 449518
rect 3969 449515 4035 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580625 418298 580691 418301
rect 583520 418298 584960 418388
rect 580625 418296 584960 418298
rect 580625 418240 580630 418296
rect 580686 418240 584960 418296
rect 580625 418238 584960 418240
rect 580625 418235 580691 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3877 358458 3943 358461
rect -960 358456 3943 358458
rect -960 358400 3882 358456
rect 3938 358400 3943 358456
rect -960 358398 3943 358400
rect -960 358308 480 358398
rect 3877 358395 3943 358398
rect 580533 351930 580599 351933
rect 583520 351930 584960 352020
rect 580533 351928 584960 351930
rect 580533 351872 580538 351928
rect 580594 351872 584960 351928
rect 580533 351870 584960 351872
rect 580533 351867 580599 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2957 345402 3023 345405
rect -960 345400 3023 345402
rect -960 345344 2962 345400
rect 3018 345344 3023 345400
rect -960 345342 3023 345344
rect -960 345252 480 345342
rect 2957 345339 3023 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 579705 312082 579771 312085
rect 583520 312082 584960 312172
rect 579705 312080 584960 312082
rect 579705 312024 579710 312080
rect 579766 312024 584960 312080
rect 579705 312022 584960 312024
rect 579705 312019 579771 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3785 306234 3851 306237
rect -960 306232 3851 306234
rect -960 306176 3790 306232
rect 3846 306176 3851 306232
rect -960 306174 3851 306176
rect -960 306084 480 306174
rect 3785 306171 3851 306174
rect 579797 298754 579863 298757
rect 583520 298754 584960 298844
rect 579797 298752 584960 298754
rect 579797 298696 579802 298752
rect 579858 298696 584960 298752
rect 579797 298694 584960 298696
rect 579797 298691 579863 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3601 241090 3667 241093
rect -960 241088 3667 241090
rect -960 241032 3606 241088
rect 3662 241032 3667 241088
rect -960 241030 3667 241032
rect -960 240940 480 241030
rect 3601 241027 3667 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 580257 192538 580323 192541
rect 583520 192538 584960 192628
rect 580257 192536 584960 192538
rect 580257 192480 580262 192536
rect 580318 192480 584960 192536
rect 580257 192478 584960 192480
rect 580257 192475 580323 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 580390 152628 580396 152692
rect 580460 152690 580466 152692
rect 583520 152690 584960 152780
rect 580460 152630 584960 152690
rect 580460 152628 580466 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 580206 139300 580212 139364
rect 580276 139362 580282 139364
rect 583520 139362 584960 139452
rect 580276 139302 584960 139362
rect 580276 139300 580282 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3734 136778 3740 136780
rect -960 136718 3740 136778
rect -960 136628 480 136718
rect 3734 136716 3740 136718
rect 3804 136716 3810 136780
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3550 84690 3556 84692
rect -960 84630 3556 84690
rect -960 84540 480 84630
rect 3550 84628 3556 84630
rect 3620 84628 3626 84692
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 579981 59666 580047 59669
rect 583520 59666 584960 59756
rect 579981 59664 584960 59666
rect 579981 59608 579986 59664
rect 580042 59608 584960 59664
rect 579981 59606 584960 59608
rect 579981 59603 580047 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3366 45522 3372 45524
rect -960 45462 3372 45522
rect -960 45372 480 45462
rect 3366 45460 3372 45462
rect 3436 45460 3442 45524
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 579797 19818 579863 19821
rect 583520 19818 584960 19908
rect 579797 19816 584960 19818
rect 579797 19760 579802 19816
rect 579858 19760 584960 19816
rect 579797 19758 584960 19760
rect 579797 19755 579863 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 579705 6626 579771 6629
rect 583520 6626 584960 6716
rect 579705 6624 584960 6626
rect -960 6490 480 6580
rect 579705 6568 579710 6624
rect 579766 6568 584960 6624
rect 579705 6566 584960 6568
rect 579705 6563 579771 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 3556 633932 3620 633996
rect 3372 633660 3436 633724
rect 580212 632300 580276 632364
rect 3740 632164 3804 632228
rect 580396 632028 580460 632092
rect 108252 631348 108316 631412
rect 108252 630668 108316 630732
rect 580396 152628 580460 152692
rect 580212 139300 580276 139364
rect 3740 136716 3804 136780
rect 3556 84628 3620 84692
rect 3372 45460 3436 45524
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 3555 633996 3621 633997
rect 3555 633932 3556 633996
rect 3620 633932 3621 633996
rect 3555 633931 3621 633932
rect 3371 633724 3437 633725
rect 3371 633660 3372 633724
rect 3436 633660 3437 633724
rect 3371 633659 3437 633660
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 45525 3434 633659
rect 3558 84693 3618 633931
rect 3739 632228 3805 632229
rect 3739 632164 3740 632228
rect 3804 632164 3805 632228
rect 3739 632163 3805 632164
rect 3742 136781 3802 632163
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 3739 136780 3805 136781
rect 3739 136716 3740 136780
rect 3804 136716 3805 136780
rect 3739 136715 3805 136716
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 3555 84692 3621 84693
rect 3555 84628 3556 84692
rect 3620 84628 3621 84692
rect 3555 84627 3621 84628
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 3371 45524 3437 45525
rect 3371 45460 3372 45524
rect 3436 45460 3437 45524
rect 3371 45459 3437 45460
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 634000 74414 650898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 634000 78914 655398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 634000 83414 659898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 634000 87914 664398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 634000 92414 668898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 634000 96914 637398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 634000 101414 641898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 634000 105914 646398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 634000 110414 650898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 634000 114914 655398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 634000 119414 659898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 634000 123914 664398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 634000 128414 668898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 634000 132914 637398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 634000 137414 641898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 634000 141914 646398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 634000 146414 650898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 634000 150914 655398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 634000 155414 659898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 634000 159914 664398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 634000 164414 668898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 634000 168914 637398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 634000 173414 641898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 634000 177914 646398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 634000 182414 650898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 634000 186914 655398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 634000 191414 659898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 634000 195914 664398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 634000 200414 668898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 634000 204914 637398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 634000 209414 641898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 634000 213914 646398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 634000 218414 650898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 634000 222914 655398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 634000 227414 659898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 634000 231914 664398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 634000 236414 668898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 634000 240914 637398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 634000 245414 641898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 634000 249914 646398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 634000 254414 650898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 634000 258914 655398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 634000 263414 659898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 634000 267914 664398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 634000 272414 668898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 634000 276914 637398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 634000 281414 641898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 634000 285914 646398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 634000 290414 650898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 634000 294914 655398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 634000 299414 659898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 634000 303914 664398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 634000 308414 668898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 634000 312914 637398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 634000 317414 641898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 634000 321914 646398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 634000 326414 650898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 634000 330914 655398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 634000 335414 659898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 634000 339914 664398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 634000 344414 668898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 634000 348914 637398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 634000 353414 641898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 634000 357914 646398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 634000 362414 650898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 634000 366914 655398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 634000 371414 659898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 634000 375914 664398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 634000 380414 668898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 634000 384914 637398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 634000 389414 641898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 634000 393914 646398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 634000 398414 650898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 634000 402914 655398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 634000 407414 659898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 634000 411914 664398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 634000 416414 668898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 634000 420914 637398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 634000 425414 641898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 634000 429914 646398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 634000 434414 650898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 634000 438914 655398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 634000 443414 659898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 634000 447914 664398
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 634000 452414 668898
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 634000 456914 637398
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 634000 461414 641898
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 634000 465914 646398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 634000 470414 650898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 634000 474914 655398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 634000 479414 659898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 634000 483914 664398
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 634000 488414 668898
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 634000 492914 637398
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 634000 497414 641898
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 634000 501914 646398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 634000 506414 650898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 634000 510914 655398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 108251 631412 108317 631413
rect 108251 631348 108252 631412
rect 108316 631348 108317 631412
rect 108251 631347 108317 631348
rect 108254 630733 108314 631347
rect 108251 630732 108317 630733
rect 108251 630668 108252 630732
rect 108316 630668 108317 630732
rect 108251 630667 108317 630668
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 91568 619954 91888 619986
rect 91568 619718 91610 619954
rect 91846 619718 91888 619954
rect 91568 619634 91888 619718
rect 91568 619398 91610 619634
rect 91846 619398 91888 619634
rect 91568 619366 91888 619398
rect 122288 619954 122608 619986
rect 122288 619718 122330 619954
rect 122566 619718 122608 619954
rect 122288 619634 122608 619718
rect 122288 619398 122330 619634
rect 122566 619398 122608 619634
rect 122288 619366 122608 619398
rect 153008 619954 153328 619986
rect 153008 619718 153050 619954
rect 153286 619718 153328 619954
rect 153008 619634 153328 619718
rect 153008 619398 153050 619634
rect 153286 619398 153328 619634
rect 153008 619366 153328 619398
rect 183728 619954 184048 619986
rect 183728 619718 183770 619954
rect 184006 619718 184048 619954
rect 183728 619634 184048 619718
rect 183728 619398 183770 619634
rect 184006 619398 184048 619634
rect 183728 619366 184048 619398
rect 214448 619954 214768 619986
rect 214448 619718 214490 619954
rect 214726 619718 214768 619954
rect 214448 619634 214768 619718
rect 214448 619398 214490 619634
rect 214726 619398 214768 619634
rect 214448 619366 214768 619398
rect 245168 619954 245488 619986
rect 245168 619718 245210 619954
rect 245446 619718 245488 619954
rect 245168 619634 245488 619718
rect 245168 619398 245210 619634
rect 245446 619398 245488 619634
rect 245168 619366 245488 619398
rect 275888 619954 276208 619986
rect 275888 619718 275930 619954
rect 276166 619718 276208 619954
rect 275888 619634 276208 619718
rect 275888 619398 275930 619634
rect 276166 619398 276208 619634
rect 275888 619366 276208 619398
rect 306608 619954 306928 619986
rect 306608 619718 306650 619954
rect 306886 619718 306928 619954
rect 306608 619634 306928 619718
rect 306608 619398 306650 619634
rect 306886 619398 306928 619634
rect 306608 619366 306928 619398
rect 337328 619954 337648 619986
rect 337328 619718 337370 619954
rect 337606 619718 337648 619954
rect 337328 619634 337648 619718
rect 337328 619398 337370 619634
rect 337606 619398 337648 619634
rect 337328 619366 337648 619398
rect 368048 619954 368368 619986
rect 368048 619718 368090 619954
rect 368326 619718 368368 619954
rect 368048 619634 368368 619718
rect 368048 619398 368090 619634
rect 368326 619398 368368 619634
rect 368048 619366 368368 619398
rect 398768 619954 399088 619986
rect 398768 619718 398810 619954
rect 399046 619718 399088 619954
rect 398768 619634 399088 619718
rect 398768 619398 398810 619634
rect 399046 619398 399088 619634
rect 398768 619366 399088 619398
rect 429488 619954 429808 619986
rect 429488 619718 429530 619954
rect 429766 619718 429808 619954
rect 429488 619634 429808 619718
rect 429488 619398 429530 619634
rect 429766 619398 429808 619634
rect 429488 619366 429808 619398
rect 460208 619954 460528 619986
rect 460208 619718 460250 619954
rect 460486 619718 460528 619954
rect 460208 619634 460528 619718
rect 460208 619398 460250 619634
rect 460486 619398 460528 619634
rect 460208 619366 460528 619398
rect 490928 619954 491248 619986
rect 490928 619718 490970 619954
rect 491206 619718 491248 619954
rect 490928 619634 491248 619718
rect 490928 619398 490970 619634
rect 491206 619398 491248 619634
rect 490928 619366 491248 619398
rect 76208 615454 76528 615486
rect 76208 615218 76250 615454
rect 76486 615218 76528 615454
rect 76208 615134 76528 615218
rect 76208 614898 76250 615134
rect 76486 614898 76528 615134
rect 76208 614866 76528 614898
rect 106928 615454 107248 615486
rect 106928 615218 106970 615454
rect 107206 615218 107248 615454
rect 106928 615134 107248 615218
rect 106928 614898 106970 615134
rect 107206 614898 107248 615134
rect 106928 614866 107248 614898
rect 137648 615454 137968 615486
rect 137648 615218 137690 615454
rect 137926 615218 137968 615454
rect 137648 615134 137968 615218
rect 137648 614898 137690 615134
rect 137926 614898 137968 615134
rect 137648 614866 137968 614898
rect 168368 615454 168688 615486
rect 168368 615218 168410 615454
rect 168646 615218 168688 615454
rect 168368 615134 168688 615218
rect 168368 614898 168410 615134
rect 168646 614898 168688 615134
rect 168368 614866 168688 614898
rect 199088 615454 199408 615486
rect 199088 615218 199130 615454
rect 199366 615218 199408 615454
rect 199088 615134 199408 615218
rect 199088 614898 199130 615134
rect 199366 614898 199408 615134
rect 199088 614866 199408 614898
rect 229808 615454 230128 615486
rect 229808 615218 229850 615454
rect 230086 615218 230128 615454
rect 229808 615134 230128 615218
rect 229808 614898 229850 615134
rect 230086 614898 230128 615134
rect 229808 614866 230128 614898
rect 260528 615454 260848 615486
rect 260528 615218 260570 615454
rect 260806 615218 260848 615454
rect 260528 615134 260848 615218
rect 260528 614898 260570 615134
rect 260806 614898 260848 615134
rect 260528 614866 260848 614898
rect 291248 615454 291568 615486
rect 291248 615218 291290 615454
rect 291526 615218 291568 615454
rect 291248 615134 291568 615218
rect 291248 614898 291290 615134
rect 291526 614898 291568 615134
rect 291248 614866 291568 614898
rect 321968 615454 322288 615486
rect 321968 615218 322010 615454
rect 322246 615218 322288 615454
rect 321968 615134 322288 615218
rect 321968 614898 322010 615134
rect 322246 614898 322288 615134
rect 321968 614866 322288 614898
rect 352688 615454 353008 615486
rect 352688 615218 352730 615454
rect 352966 615218 353008 615454
rect 352688 615134 353008 615218
rect 352688 614898 352730 615134
rect 352966 614898 353008 615134
rect 352688 614866 353008 614898
rect 383408 615454 383728 615486
rect 383408 615218 383450 615454
rect 383686 615218 383728 615454
rect 383408 615134 383728 615218
rect 383408 614898 383450 615134
rect 383686 614898 383728 615134
rect 383408 614866 383728 614898
rect 414128 615454 414448 615486
rect 414128 615218 414170 615454
rect 414406 615218 414448 615454
rect 414128 615134 414448 615218
rect 414128 614898 414170 615134
rect 414406 614898 414448 615134
rect 414128 614866 414448 614898
rect 444848 615454 445168 615486
rect 444848 615218 444890 615454
rect 445126 615218 445168 615454
rect 444848 615134 445168 615218
rect 444848 614898 444890 615134
rect 445126 614898 445168 615134
rect 444848 614866 445168 614898
rect 475568 615454 475888 615486
rect 475568 615218 475610 615454
rect 475846 615218 475888 615454
rect 475568 615134 475888 615218
rect 475568 614898 475610 615134
rect 475846 614898 475888 615134
rect 475568 614866 475888 614898
rect 506288 615454 506608 615486
rect 506288 615218 506330 615454
rect 506566 615218 506608 615454
rect 506288 615134 506608 615218
rect 506288 614898 506330 615134
rect 506566 614898 506608 615134
rect 506288 614866 506608 614898
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 91568 583954 91888 583986
rect 91568 583718 91610 583954
rect 91846 583718 91888 583954
rect 91568 583634 91888 583718
rect 91568 583398 91610 583634
rect 91846 583398 91888 583634
rect 91568 583366 91888 583398
rect 122288 583954 122608 583986
rect 122288 583718 122330 583954
rect 122566 583718 122608 583954
rect 122288 583634 122608 583718
rect 122288 583398 122330 583634
rect 122566 583398 122608 583634
rect 122288 583366 122608 583398
rect 153008 583954 153328 583986
rect 153008 583718 153050 583954
rect 153286 583718 153328 583954
rect 153008 583634 153328 583718
rect 153008 583398 153050 583634
rect 153286 583398 153328 583634
rect 153008 583366 153328 583398
rect 183728 583954 184048 583986
rect 183728 583718 183770 583954
rect 184006 583718 184048 583954
rect 183728 583634 184048 583718
rect 183728 583398 183770 583634
rect 184006 583398 184048 583634
rect 183728 583366 184048 583398
rect 214448 583954 214768 583986
rect 214448 583718 214490 583954
rect 214726 583718 214768 583954
rect 214448 583634 214768 583718
rect 214448 583398 214490 583634
rect 214726 583398 214768 583634
rect 214448 583366 214768 583398
rect 245168 583954 245488 583986
rect 245168 583718 245210 583954
rect 245446 583718 245488 583954
rect 245168 583634 245488 583718
rect 245168 583398 245210 583634
rect 245446 583398 245488 583634
rect 245168 583366 245488 583398
rect 275888 583954 276208 583986
rect 275888 583718 275930 583954
rect 276166 583718 276208 583954
rect 275888 583634 276208 583718
rect 275888 583398 275930 583634
rect 276166 583398 276208 583634
rect 275888 583366 276208 583398
rect 306608 583954 306928 583986
rect 306608 583718 306650 583954
rect 306886 583718 306928 583954
rect 306608 583634 306928 583718
rect 306608 583398 306650 583634
rect 306886 583398 306928 583634
rect 306608 583366 306928 583398
rect 337328 583954 337648 583986
rect 337328 583718 337370 583954
rect 337606 583718 337648 583954
rect 337328 583634 337648 583718
rect 337328 583398 337370 583634
rect 337606 583398 337648 583634
rect 337328 583366 337648 583398
rect 368048 583954 368368 583986
rect 368048 583718 368090 583954
rect 368326 583718 368368 583954
rect 368048 583634 368368 583718
rect 368048 583398 368090 583634
rect 368326 583398 368368 583634
rect 368048 583366 368368 583398
rect 398768 583954 399088 583986
rect 398768 583718 398810 583954
rect 399046 583718 399088 583954
rect 398768 583634 399088 583718
rect 398768 583398 398810 583634
rect 399046 583398 399088 583634
rect 398768 583366 399088 583398
rect 429488 583954 429808 583986
rect 429488 583718 429530 583954
rect 429766 583718 429808 583954
rect 429488 583634 429808 583718
rect 429488 583398 429530 583634
rect 429766 583398 429808 583634
rect 429488 583366 429808 583398
rect 460208 583954 460528 583986
rect 460208 583718 460250 583954
rect 460486 583718 460528 583954
rect 460208 583634 460528 583718
rect 460208 583398 460250 583634
rect 460486 583398 460528 583634
rect 460208 583366 460528 583398
rect 490928 583954 491248 583986
rect 490928 583718 490970 583954
rect 491206 583718 491248 583954
rect 490928 583634 491248 583718
rect 490928 583398 490970 583634
rect 491206 583398 491248 583634
rect 490928 583366 491248 583398
rect 76208 579454 76528 579486
rect 76208 579218 76250 579454
rect 76486 579218 76528 579454
rect 76208 579134 76528 579218
rect 76208 578898 76250 579134
rect 76486 578898 76528 579134
rect 76208 578866 76528 578898
rect 106928 579454 107248 579486
rect 106928 579218 106970 579454
rect 107206 579218 107248 579454
rect 106928 579134 107248 579218
rect 106928 578898 106970 579134
rect 107206 578898 107248 579134
rect 106928 578866 107248 578898
rect 137648 579454 137968 579486
rect 137648 579218 137690 579454
rect 137926 579218 137968 579454
rect 137648 579134 137968 579218
rect 137648 578898 137690 579134
rect 137926 578898 137968 579134
rect 137648 578866 137968 578898
rect 168368 579454 168688 579486
rect 168368 579218 168410 579454
rect 168646 579218 168688 579454
rect 168368 579134 168688 579218
rect 168368 578898 168410 579134
rect 168646 578898 168688 579134
rect 168368 578866 168688 578898
rect 199088 579454 199408 579486
rect 199088 579218 199130 579454
rect 199366 579218 199408 579454
rect 199088 579134 199408 579218
rect 199088 578898 199130 579134
rect 199366 578898 199408 579134
rect 199088 578866 199408 578898
rect 229808 579454 230128 579486
rect 229808 579218 229850 579454
rect 230086 579218 230128 579454
rect 229808 579134 230128 579218
rect 229808 578898 229850 579134
rect 230086 578898 230128 579134
rect 229808 578866 230128 578898
rect 260528 579454 260848 579486
rect 260528 579218 260570 579454
rect 260806 579218 260848 579454
rect 260528 579134 260848 579218
rect 260528 578898 260570 579134
rect 260806 578898 260848 579134
rect 260528 578866 260848 578898
rect 291248 579454 291568 579486
rect 291248 579218 291290 579454
rect 291526 579218 291568 579454
rect 291248 579134 291568 579218
rect 291248 578898 291290 579134
rect 291526 578898 291568 579134
rect 291248 578866 291568 578898
rect 321968 579454 322288 579486
rect 321968 579218 322010 579454
rect 322246 579218 322288 579454
rect 321968 579134 322288 579218
rect 321968 578898 322010 579134
rect 322246 578898 322288 579134
rect 321968 578866 322288 578898
rect 352688 579454 353008 579486
rect 352688 579218 352730 579454
rect 352966 579218 353008 579454
rect 352688 579134 353008 579218
rect 352688 578898 352730 579134
rect 352966 578898 353008 579134
rect 352688 578866 353008 578898
rect 383408 579454 383728 579486
rect 383408 579218 383450 579454
rect 383686 579218 383728 579454
rect 383408 579134 383728 579218
rect 383408 578898 383450 579134
rect 383686 578898 383728 579134
rect 383408 578866 383728 578898
rect 414128 579454 414448 579486
rect 414128 579218 414170 579454
rect 414406 579218 414448 579454
rect 414128 579134 414448 579218
rect 414128 578898 414170 579134
rect 414406 578898 414448 579134
rect 414128 578866 414448 578898
rect 444848 579454 445168 579486
rect 444848 579218 444890 579454
rect 445126 579218 445168 579454
rect 444848 579134 445168 579218
rect 444848 578898 444890 579134
rect 445126 578898 445168 579134
rect 444848 578866 445168 578898
rect 475568 579454 475888 579486
rect 475568 579218 475610 579454
rect 475846 579218 475888 579454
rect 475568 579134 475888 579218
rect 475568 578898 475610 579134
rect 475846 578898 475888 579134
rect 475568 578866 475888 578898
rect 506288 579454 506608 579486
rect 506288 579218 506330 579454
rect 506566 579218 506608 579454
rect 506288 579134 506608 579218
rect 506288 578898 506330 579134
rect 506566 578898 506608 579134
rect 506288 578866 506608 578898
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 91568 547954 91888 547986
rect 91568 547718 91610 547954
rect 91846 547718 91888 547954
rect 91568 547634 91888 547718
rect 91568 547398 91610 547634
rect 91846 547398 91888 547634
rect 91568 547366 91888 547398
rect 122288 547954 122608 547986
rect 122288 547718 122330 547954
rect 122566 547718 122608 547954
rect 122288 547634 122608 547718
rect 122288 547398 122330 547634
rect 122566 547398 122608 547634
rect 122288 547366 122608 547398
rect 153008 547954 153328 547986
rect 153008 547718 153050 547954
rect 153286 547718 153328 547954
rect 153008 547634 153328 547718
rect 153008 547398 153050 547634
rect 153286 547398 153328 547634
rect 153008 547366 153328 547398
rect 183728 547954 184048 547986
rect 183728 547718 183770 547954
rect 184006 547718 184048 547954
rect 183728 547634 184048 547718
rect 183728 547398 183770 547634
rect 184006 547398 184048 547634
rect 183728 547366 184048 547398
rect 214448 547954 214768 547986
rect 214448 547718 214490 547954
rect 214726 547718 214768 547954
rect 214448 547634 214768 547718
rect 214448 547398 214490 547634
rect 214726 547398 214768 547634
rect 214448 547366 214768 547398
rect 245168 547954 245488 547986
rect 245168 547718 245210 547954
rect 245446 547718 245488 547954
rect 245168 547634 245488 547718
rect 245168 547398 245210 547634
rect 245446 547398 245488 547634
rect 245168 547366 245488 547398
rect 275888 547954 276208 547986
rect 275888 547718 275930 547954
rect 276166 547718 276208 547954
rect 275888 547634 276208 547718
rect 275888 547398 275930 547634
rect 276166 547398 276208 547634
rect 275888 547366 276208 547398
rect 306608 547954 306928 547986
rect 306608 547718 306650 547954
rect 306886 547718 306928 547954
rect 306608 547634 306928 547718
rect 306608 547398 306650 547634
rect 306886 547398 306928 547634
rect 306608 547366 306928 547398
rect 337328 547954 337648 547986
rect 337328 547718 337370 547954
rect 337606 547718 337648 547954
rect 337328 547634 337648 547718
rect 337328 547398 337370 547634
rect 337606 547398 337648 547634
rect 337328 547366 337648 547398
rect 368048 547954 368368 547986
rect 368048 547718 368090 547954
rect 368326 547718 368368 547954
rect 368048 547634 368368 547718
rect 368048 547398 368090 547634
rect 368326 547398 368368 547634
rect 368048 547366 368368 547398
rect 398768 547954 399088 547986
rect 398768 547718 398810 547954
rect 399046 547718 399088 547954
rect 398768 547634 399088 547718
rect 398768 547398 398810 547634
rect 399046 547398 399088 547634
rect 398768 547366 399088 547398
rect 429488 547954 429808 547986
rect 429488 547718 429530 547954
rect 429766 547718 429808 547954
rect 429488 547634 429808 547718
rect 429488 547398 429530 547634
rect 429766 547398 429808 547634
rect 429488 547366 429808 547398
rect 460208 547954 460528 547986
rect 460208 547718 460250 547954
rect 460486 547718 460528 547954
rect 460208 547634 460528 547718
rect 460208 547398 460250 547634
rect 460486 547398 460528 547634
rect 460208 547366 460528 547398
rect 490928 547954 491248 547986
rect 490928 547718 490970 547954
rect 491206 547718 491248 547954
rect 490928 547634 491248 547718
rect 490928 547398 490970 547634
rect 491206 547398 491248 547634
rect 490928 547366 491248 547398
rect 76208 543454 76528 543486
rect 76208 543218 76250 543454
rect 76486 543218 76528 543454
rect 76208 543134 76528 543218
rect 76208 542898 76250 543134
rect 76486 542898 76528 543134
rect 76208 542866 76528 542898
rect 106928 543454 107248 543486
rect 106928 543218 106970 543454
rect 107206 543218 107248 543454
rect 106928 543134 107248 543218
rect 106928 542898 106970 543134
rect 107206 542898 107248 543134
rect 106928 542866 107248 542898
rect 137648 543454 137968 543486
rect 137648 543218 137690 543454
rect 137926 543218 137968 543454
rect 137648 543134 137968 543218
rect 137648 542898 137690 543134
rect 137926 542898 137968 543134
rect 137648 542866 137968 542898
rect 168368 543454 168688 543486
rect 168368 543218 168410 543454
rect 168646 543218 168688 543454
rect 168368 543134 168688 543218
rect 168368 542898 168410 543134
rect 168646 542898 168688 543134
rect 168368 542866 168688 542898
rect 199088 543454 199408 543486
rect 199088 543218 199130 543454
rect 199366 543218 199408 543454
rect 199088 543134 199408 543218
rect 199088 542898 199130 543134
rect 199366 542898 199408 543134
rect 199088 542866 199408 542898
rect 229808 543454 230128 543486
rect 229808 543218 229850 543454
rect 230086 543218 230128 543454
rect 229808 543134 230128 543218
rect 229808 542898 229850 543134
rect 230086 542898 230128 543134
rect 229808 542866 230128 542898
rect 260528 543454 260848 543486
rect 260528 543218 260570 543454
rect 260806 543218 260848 543454
rect 260528 543134 260848 543218
rect 260528 542898 260570 543134
rect 260806 542898 260848 543134
rect 260528 542866 260848 542898
rect 291248 543454 291568 543486
rect 291248 543218 291290 543454
rect 291526 543218 291568 543454
rect 291248 543134 291568 543218
rect 291248 542898 291290 543134
rect 291526 542898 291568 543134
rect 291248 542866 291568 542898
rect 321968 543454 322288 543486
rect 321968 543218 322010 543454
rect 322246 543218 322288 543454
rect 321968 543134 322288 543218
rect 321968 542898 322010 543134
rect 322246 542898 322288 543134
rect 321968 542866 322288 542898
rect 352688 543454 353008 543486
rect 352688 543218 352730 543454
rect 352966 543218 353008 543454
rect 352688 543134 353008 543218
rect 352688 542898 352730 543134
rect 352966 542898 353008 543134
rect 352688 542866 353008 542898
rect 383408 543454 383728 543486
rect 383408 543218 383450 543454
rect 383686 543218 383728 543454
rect 383408 543134 383728 543218
rect 383408 542898 383450 543134
rect 383686 542898 383728 543134
rect 383408 542866 383728 542898
rect 414128 543454 414448 543486
rect 414128 543218 414170 543454
rect 414406 543218 414448 543454
rect 414128 543134 414448 543218
rect 414128 542898 414170 543134
rect 414406 542898 414448 543134
rect 414128 542866 414448 542898
rect 444848 543454 445168 543486
rect 444848 543218 444890 543454
rect 445126 543218 445168 543454
rect 444848 543134 445168 543218
rect 444848 542898 444890 543134
rect 445126 542898 445168 543134
rect 444848 542866 445168 542898
rect 475568 543454 475888 543486
rect 475568 543218 475610 543454
rect 475846 543218 475888 543454
rect 475568 543134 475888 543218
rect 475568 542898 475610 543134
rect 475846 542898 475888 543134
rect 475568 542866 475888 542898
rect 506288 543454 506608 543486
rect 506288 543218 506330 543454
rect 506566 543218 506608 543454
rect 506288 543134 506608 543218
rect 506288 542898 506330 543134
rect 506566 542898 506608 543134
rect 506288 542866 506608 542898
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 91568 511954 91888 511986
rect 91568 511718 91610 511954
rect 91846 511718 91888 511954
rect 91568 511634 91888 511718
rect 91568 511398 91610 511634
rect 91846 511398 91888 511634
rect 91568 511366 91888 511398
rect 122288 511954 122608 511986
rect 122288 511718 122330 511954
rect 122566 511718 122608 511954
rect 122288 511634 122608 511718
rect 122288 511398 122330 511634
rect 122566 511398 122608 511634
rect 122288 511366 122608 511398
rect 153008 511954 153328 511986
rect 153008 511718 153050 511954
rect 153286 511718 153328 511954
rect 153008 511634 153328 511718
rect 153008 511398 153050 511634
rect 153286 511398 153328 511634
rect 153008 511366 153328 511398
rect 183728 511954 184048 511986
rect 183728 511718 183770 511954
rect 184006 511718 184048 511954
rect 183728 511634 184048 511718
rect 183728 511398 183770 511634
rect 184006 511398 184048 511634
rect 183728 511366 184048 511398
rect 214448 511954 214768 511986
rect 214448 511718 214490 511954
rect 214726 511718 214768 511954
rect 214448 511634 214768 511718
rect 214448 511398 214490 511634
rect 214726 511398 214768 511634
rect 214448 511366 214768 511398
rect 245168 511954 245488 511986
rect 245168 511718 245210 511954
rect 245446 511718 245488 511954
rect 245168 511634 245488 511718
rect 245168 511398 245210 511634
rect 245446 511398 245488 511634
rect 245168 511366 245488 511398
rect 275888 511954 276208 511986
rect 275888 511718 275930 511954
rect 276166 511718 276208 511954
rect 275888 511634 276208 511718
rect 275888 511398 275930 511634
rect 276166 511398 276208 511634
rect 275888 511366 276208 511398
rect 306608 511954 306928 511986
rect 306608 511718 306650 511954
rect 306886 511718 306928 511954
rect 306608 511634 306928 511718
rect 306608 511398 306650 511634
rect 306886 511398 306928 511634
rect 306608 511366 306928 511398
rect 337328 511954 337648 511986
rect 337328 511718 337370 511954
rect 337606 511718 337648 511954
rect 337328 511634 337648 511718
rect 337328 511398 337370 511634
rect 337606 511398 337648 511634
rect 337328 511366 337648 511398
rect 368048 511954 368368 511986
rect 368048 511718 368090 511954
rect 368326 511718 368368 511954
rect 368048 511634 368368 511718
rect 368048 511398 368090 511634
rect 368326 511398 368368 511634
rect 368048 511366 368368 511398
rect 398768 511954 399088 511986
rect 398768 511718 398810 511954
rect 399046 511718 399088 511954
rect 398768 511634 399088 511718
rect 398768 511398 398810 511634
rect 399046 511398 399088 511634
rect 398768 511366 399088 511398
rect 429488 511954 429808 511986
rect 429488 511718 429530 511954
rect 429766 511718 429808 511954
rect 429488 511634 429808 511718
rect 429488 511398 429530 511634
rect 429766 511398 429808 511634
rect 429488 511366 429808 511398
rect 460208 511954 460528 511986
rect 460208 511718 460250 511954
rect 460486 511718 460528 511954
rect 460208 511634 460528 511718
rect 460208 511398 460250 511634
rect 460486 511398 460528 511634
rect 460208 511366 460528 511398
rect 490928 511954 491248 511986
rect 490928 511718 490970 511954
rect 491206 511718 491248 511954
rect 490928 511634 491248 511718
rect 490928 511398 490970 511634
rect 491206 511398 491248 511634
rect 490928 511366 491248 511398
rect 76208 507454 76528 507486
rect 76208 507218 76250 507454
rect 76486 507218 76528 507454
rect 76208 507134 76528 507218
rect 76208 506898 76250 507134
rect 76486 506898 76528 507134
rect 76208 506866 76528 506898
rect 106928 507454 107248 507486
rect 106928 507218 106970 507454
rect 107206 507218 107248 507454
rect 106928 507134 107248 507218
rect 106928 506898 106970 507134
rect 107206 506898 107248 507134
rect 106928 506866 107248 506898
rect 137648 507454 137968 507486
rect 137648 507218 137690 507454
rect 137926 507218 137968 507454
rect 137648 507134 137968 507218
rect 137648 506898 137690 507134
rect 137926 506898 137968 507134
rect 137648 506866 137968 506898
rect 168368 507454 168688 507486
rect 168368 507218 168410 507454
rect 168646 507218 168688 507454
rect 168368 507134 168688 507218
rect 168368 506898 168410 507134
rect 168646 506898 168688 507134
rect 168368 506866 168688 506898
rect 199088 507454 199408 507486
rect 199088 507218 199130 507454
rect 199366 507218 199408 507454
rect 199088 507134 199408 507218
rect 199088 506898 199130 507134
rect 199366 506898 199408 507134
rect 199088 506866 199408 506898
rect 229808 507454 230128 507486
rect 229808 507218 229850 507454
rect 230086 507218 230128 507454
rect 229808 507134 230128 507218
rect 229808 506898 229850 507134
rect 230086 506898 230128 507134
rect 229808 506866 230128 506898
rect 260528 507454 260848 507486
rect 260528 507218 260570 507454
rect 260806 507218 260848 507454
rect 260528 507134 260848 507218
rect 260528 506898 260570 507134
rect 260806 506898 260848 507134
rect 260528 506866 260848 506898
rect 291248 507454 291568 507486
rect 291248 507218 291290 507454
rect 291526 507218 291568 507454
rect 291248 507134 291568 507218
rect 291248 506898 291290 507134
rect 291526 506898 291568 507134
rect 291248 506866 291568 506898
rect 321968 507454 322288 507486
rect 321968 507218 322010 507454
rect 322246 507218 322288 507454
rect 321968 507134 322288 507218
rect 321968 506898 322010 507134
rect 322246 506898 322288 507134
rect 321968 506866 322288 506898
rect 352688 507454 353008 507486
rect 352688 507218 352730 507454
rect 352966 507218 353008 507454
rect 352688 507134 353008 507218
rect 352688 506898 352730 507134
rect 352966 506898 353008 507134
rect 352688 506866 353008 506898
rect 383408 507454 383728 507486
rect 383408 507218 383450 507454
rect 383686 507218 383728 507454
rect 383408 507134 383728 507218
rect 383408 506898 383450 507134
rect 383686 506898 383728 507134
rect 383408 506866 383728 506898
rect 414128 507454 414448 507486
rect 414128 507218 414170 507454
rect 414406 507218 414448 507454
rect 414128 507134 414448 507218
rect 414128 506898 414170 507134
rect 414406 506898 414448 507134
rect 414128 506866 414448 506898
rect 444848 507454 445168 507486
rect 444848 507218 444890 507454
rect 445126 507218 445168 507454
rect 444848 507134 445168 507218
rect 444848 506898 444890 507134
rect 445126 506898 445168 507134
rect 444848 506866 445168 506898
rect 475568 507454 475888 507486
rect 475568 507218 475610 507454
rect 475846 507218 475888 507454
rect 475568 507134 475888 507218
rect 475568 506898 475610 507134
rect 475846 506898 475888 507134
rect 475568 506866 475888 506898
rect 506288 507454 506608 507486
rect 506288 507218 506330 507454
rect 506566 507218 506608 507454
rect 506288 507134 506608 507218
rect 506288 506898 506330 507134
rect 506566 506898 506608 507134
rect 506288 506866 506608 506898
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 91568 475954 91888 475986
rect 91568 475718 91610 475954
rect 91846 475718 91888 475954
rect 91568 475634 91888 475718
rect 91568 475398 91610 475634
rect 91846 475398 91888 475634
rect 91568 475366 91888 475398
rect 122288 475954 122608 475986
rect 122288 475718 122330 475954
rect 122566 475718 122608 475954
rect 122288 475634 122608 475718
rect 122288 475398 122330 475634
rect 122566 475398 122608 475634
rect 122288 475366 122608 475398
rect 153008 475954 153328 475986
rect 153008 475718 153050 475954
rect 153286 475718 153328 475954
rect 153008 475634 153328 475718
rect 153008 475398 153050 475634
rect 153286 475398 153328 475634
rect 153008 475366 153328 475398
rect 183728 475954 184048 475986
rect 183728 475718 183770 475954
rect 184006 475718 184048 475954
rect 183728 475634 184048 475718
rect 183728 475398 183770 475634
rect 184006 475398 184048 475634
rect 183728 475366 184048 475398
rect 214448 475954 214768 475986
rect 214448 475718 214490 475954
rect 214726 475718 214768 475954
rect 214448 475634 214768 475718
rect 214448 475398 214490 475634
rect 214726 475398 214768 475634
rect 214448 475366 214768 475398
rect 245168 475954 245488 475986
rect 245168 475718 245210 475954
rect 245446 475718 245488 475954
rect 245168 475634 245488 475718
rect 245168 475398 245210 475634
rect 245446 475398 245488 475634
rect 245168 475366 245488 475398
rect 275888 475954 276208 475986
rect 275888 475718 275930 475954
rect 276166 475718 276208 475954
rect 275888 475634 276208 475718
rect 275888 475398 275930 475634
rect 276166 475398 276208 475634
rect 275888 475366 276208 475398
rect 306608 475954 306928 475986
rect 306608 475718 306650 475954
rect 306886 475718 306928 475954
rect 306608 475634 306928 475718
rect 306608 475398 306650 475634
rect 306886 475398 306928 475634
rect 306608 475366 306928 475398
rect 337328 475954 337648 475986
rect 337328 475718 337370 475954
rect 337606 475718 337648 475954
rect 337328 475634 337648 475718
rect 337328 475398 337370 475634
rect 337606 475398 337648 475634
rect 337328 475366 337648 475398
rect 368048 475954 368368 475986
rect 368048 475718 368090 475954
rect 368326 475718 368368 475954
rect 368048 475634 368368 475718
rect 368048 475398 368090 475634
rect 368326 475398 368368 475634
rect 368048 475366 368368 475398
rect 398768 475954 399088 475986
rect 398768 475718 398810 475954
rect 399046 475718 399088 475954
rect 398768 475634 399088 475718
rect 398768 475398 398810 475634
rect 399046 475398 399088 475634
rect 398768 475366 399088 475398
rect 429488 475954 429808 475986
rect 429488 475718 429530 475954
rect 429766 475718 429808 475954
rect 429488 475634 429808 475718
rect 429488 475398 429530 475634
rect 429766 475398 429808 475634
rect 429488 475366 429808 475398
rect 460208 475954 460528 475986
rect 460208 475718 460250 475954
rect 460486 475718 460528 475954
rect 460208 475634 460528 475718
rect 460208 475398 460250 475634
rect 460486 475398 460528 475634
rect 460208 475366 460528 475398
rect 490928 475954 491248 475986
rect 490928 475718 490970 475954
rect 491206 475718 491248 475954
rect 490928 475634 491248 475718
rect 490928 475398 490970 475634
rect 491206 475398 491248 475634
rect 490928 475366 491248 475398
rect 76208 471454 76528 471486
rect 76208 471218 76250 471454
rect 76486 471218 76528 471454
rect 76208 471134 76528 471218
rect 76208 470898 76250 471134
rect 76486 470898 76528 471134
rect 76208 470866 76528 470898
rect 106928 471454 107248 471486
rect 106928 471218 106970 471454
rect 107206 471218 107248 471454
rect 106928 471134 107248 471218
rect 106928 470898 106970 471134
rect 107206 470898 107248 471134
rect 106928 470866 107248 470898
rect 137648 471454 137968 471486
rect 137648 471218 137690 471454
rect 137926 471218 137968 471454
rect 137648 471134 137968 471218
rect 137648 470898 137690 471134
rect 137926 470898 137968 471134
rect 137648 470866 137968 470898
rect 168368 471454 168688 471486
rect 168368 471218 168410 471454
rect 168646 471218 168688 471454
rect 168368 471134 168688 471218
rect 168368 470898 168410 471134
rect 168646 470898 168688 471134
rect 168368 470866 168688 470898
rect 199088 471454 199408 471486
rect 199088 471218 199130 471454
rect 199366 471218 199408 471454
rect 199088 471134 199408 471218
rect 199088 470898 199130 471134
rect 199366 470898 199408 471134
rect 199088 470866 199408 470898
rect 229808 471454 230128 471486
rect 229808 471218 229850 471454
rect 230086 471218 230128 471454
rect 229808 471134 230128 471218
rect 229808 470898 229850 471134
rect 230086 470898 230128 471134
rect 229808 470866 230128 470898
rect 260528 471454 260848 471486
rect 260528 471218 260570 471454
rect 260806 471218 260848 471454
rect 260528 471134 260848 471218
rect 260528 470898 260570 471134
rect 260806 470898 260848 471134
rect 260528 470866 260848 470898
rect 291248 471454 291568 471486
rect 291248 471218 291290 471454
rect 291526 471218 291568 471454
rect 291248 471134 291568 471218
rect 291248 470898 291290 471134
rect 291526 470898 291568 471134
rect 291248 470866 291568 470898
rect 321968 471454 322288 471486
rect 321968 471218 322010 471454
rect 322246 471218 322288 471454
rect 321968 471134 322288 471218
rect 321968 470898 322010 471134
rect 322246 470898 322288 471134
rect 321968 470866 322288 470898
rect 352688 471454 353008 471486
rect 352688 471218 352730 471454
rect 352966 471218 353008 471454
rect 352688 471134 353008 471218
rect 352688 470898 352730 471134
rect 352966 470898 353008 471134
rect 352688 470866 353008 470898
rect 383408 471454 383728 471486
rect 383408 471218 383450 471454
rect 383686 471218 383728 471454
rect 383408 471134 383728 471218
rect 383408 470898 383450 471134
rect 383686 470898 383728 471134
rect 383408 470866 383728 470898
rect 414128 471454 414448 471486
rect 414128 471218 414170 471454
rect 414406 471218 414448 471454
rect 414128 471134 414448 471218
rect 414128 470898 414170 471134
rect 414406 470898 414448 471134
rect 414128 470866 414448 470898
rect 444848 471454 445168 471486
rect 444848 471218 444890 471454
rect 445126 471218 445168 471454
rect 444848 471134 445168 471218
rect 444848 470898 444890 471134
rect 445126 470898 445168 471134
rect 444848 470866 445168 470898
rect 475568 471454 475888 471486
rect 475568 471218 475610 471454
rect 475846 471218 475888 471454
rect 475568 471134 475888 471218
rect 475568 470898 475610 471134
rect 475846 470898 475888 471134
rect 475568 470866 475888 470898
rect 506288 471454 506608 471486
rect 506288 471218 506330 471454
rect 506566 471218 506608 471454
rect 506288 471134 506608 471218
rect 506288 470898 506330 471134
rect 506566 470898 506608 471134
rect 506288 470866 506608 470898
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 91568 439954 91888 439986
rect 91568 439718 91610 439954
rect 91846 439718 91888 439954
rect 91568 439634 91888 439718
rect 91568 439398 91610 439634
rect 91846 439398 91888 439634
rect 91568 439366 91888 439398
rect 122288 439954 122608 439986
rect 122288 439718 122330 439954
rect 122566 439718 122608 439954
rect 122288 439634 122608 439718
rect 122288 439398 122330 439634
rect 122566 439398 122608 439634
rect 122288 439366 122608 439398
rect 153008 439954 153328 439986
rect 153008 439718 153050 439954
rect 153286 439718 153328 439954
rect 153008 439634 153328 439718
rect 153008 439398 153050 439634
rect 153286 439398 153328 439634
rect 153008 439366 153328 439398
rect 183728 439954 184048 439986
rect 183728 439718 183770 439954
rect 184006 439718 184048 439954
rect 183728 439634 184048 439718
rect 183728 439398 183770 439634
rect 184006 439398 184048 439634
rect 183728 439366 184048 439398
rect 214448 439954 214768 439986
rect 214448 439718 214490 439954
rect 214726 439718 214768 439954
rect 214448 439634 214768 439718
rect 214448 439398 214490 439634
rect 214726 439398 214768 439634
rect 214448 439366 214768 439398
rect 245168 439954 245488 439986
rect 245168 439718 245210 439954
rect 245446 439718 245488 439954
rect 245168 439634 245488 439718
rect 245168 439398 245210 439634
rect 245446 439398 245488 439634
rect 245168 439366 245488 439398
rect 275888 439954 276208 439986
rect 275888 439718 275930 439954
rect 276166 439718 276208 439954
rect 275888 439634 276208 439718
rect 275888 439398 275930 439634
rect 276166 439398 276208 439634
rect 275888 439366 276208 439398
rect 306608 439954 306928 439986
rect 306608 439718 306650 439954
rect 306886 439718 306928 439954
rect 306608 439634 306928 439718
rect 306608 439398 306650 439634
rect 306886 439398 306928 439634
rect 306608 439366 306928 439398
rect 337328 439954 337648 439986
rect 337328 439718 337370 439954
rect 337606 439718 337648 439954
rect 337328 439634 337648 439718
rect 337328 439398 337370 439634
rect 337606 439398 337648 439634
rect 337328 439366 337648 439398
rect 368048 439954 368368 439986
rect 368048 439718 368090 439954
rect 368326 439718 368368 439954
rect 368048 439634 368368 439718
rect 368048 439398 368090 439634
rect 368326 439398 368368 439634
rect 368048 439366 368368 439398
rect 398768 439954 399088 439986
rect 398768 439718 398810 439954
rect 399046 439718 399088 439954
rect 398768 439634 399088 439718
rect 398768 439398 398810 439634
rect 399046 439398 399088 439634
rect 398768 439366 399088 439398
rect 429488 439954 429808 439986
rect 429488 439718 429530 439954
rect 429766 439718 429808 439954
rect 429488 439634 429808 439718
rect 429488 439398 429530 439634
rect 429766 439398 429808 439634
rect 429488 439366 429808 439398
rect 460208 439954 460528 439986
rect 460208 439718 460250 439954
rect 460486 439718 460528 439954
rect 460208 439634 460528 439718
rect 460208 439398 460250 439634
rect 460486 439398 460528 439634
rect 460208 439366 460528 439398
rect 490928 439954 491248 439986
rect 490928 439718 490970 439954
rect 491206 439718 491248 439954
rect 490928 439634 491248 439718
rect 490928 439398 490970 439634
rect 491206 439398 491248 439634
rect 490928 439366 491248 439398
rect 76208 435454 76528 435486
rect 76208 435218 76250 435454
rect 76486 435218 76528 435454
rect 76208 435134 76528 435218
rect 76208 434898 76250 435134
rect 76486 434898 76528 435134
rect 76208 434866 76528 434898
rect 106928 435454 107248 435486
rect 106928 435218 106970 435454
rect 107206 435218 107248 435454
rect 106928 435134 107248 435218
rect 106928 434898 106970 435134
rect 107206 434898 107248 435134
rect 106928 434866 107248 434898
rect 137648 435454 137968 435486
rect 137648 435218 137690 435454
rect 137926 435218 137968 435454
rect 137648 435134 137968 435218
rect 137648 434898 137690 435134
rect 137926 434898 137968 435134
rect 137648 434866 137968 434898
rect 168368 435454 168688 435486
rect 168368 435218 168410 435454
rect 168646 435218 168688 435454
rect 168368 435134 168688 435218
rect 168368 434898 168410 435134
rect 168646 434898 168688 435134
rect 168368 434866 168688 434898
rect 199088 435454 199408 435486
rect 199088 435218 199130 435454
rect 199366 435218 199408 435454
rect 199088 435134 199408 435218
rect 199088 434898 199130 435134
rect 199366 434898 199408 435134
rect 199088 434866 199408 434898
rect 229808 435454 230128 435486
rect 229808 435218 229850 435454
rect 230086 435218 230128 435454
rect 229808 435134 230128 435218
rect 229808 434898 229850 435134
rect 230086 434898 230128 435134
rect 229808 434866 230128 434898
rect 260528 435454 260848 435486
rect 260528 435218 260570 435454
rect 260806 435218 260848 435454
rect 260528 435134 260848 435218
rect 260528 434898 260570 435134
rect 260806 434898 260848 435134
rect 260528 434866 260848 434898
rect 291248 435454 291568 435486
rect 291248 435218 291290 435454
rect 291526 435218 291568 435454
rect 291248 435134 291568 435218
rect 291248 434898 291290 435134
rect 291526 434898 291568 435134
rect 291248 434866 291568 434898
rect 321968 435454 322288 435486
rect 321968 435218 322010 435454
rect 322246 435218 322288 435454
rect 321968 435134 322288 435218
rect 321968 434898 322010 435134
rect 322246 434898 322288 435134
rect 321968 434866 322288 434898
rect 352688 435454 353008 435486
rect 352688 435218 352730 435454
rect 352966 435218 353008 435454
rect 352688 435134 353008 435218
rect 352688 434898 352730 435134
rect 352966 434898 353008 435134
rect 352688 434866 353008 434898
rect 383408 435454 383728 435486
rect 383408 435218 383450 435454
rect 383686 435218 383728 435454
rect 383408 435134 383728 435218
rect 383408 434898 383450 435134
rect 383686 434898 383728 435134
rect 383408 434866 383728 434898
rect 414128 435454 414448 435486
rect 414128 435218 414170 435454
rect 414406 435218 414448 435454
rect 414128 435134 414448 435218
rect 414128 434898 414170 435134
rect 414406 434898 414448 435134
rect 414128 434866 414448 434898
rect 444848 435454 445168 435486
rect 444848 435218 444890 435454
rect 445126 435218 445168 435454
rect 444848 435134 445168 435218
rect 444848 434898 444890 435134
rect 445126 434898 445168 435134
rect 444848 434866 445168 434898
rect 475568 435454 475888 435486
rect 475568 435218 475610 435454
rect 475846 435218 475888 435454
rect 475568 435134 475888 435218
rect 475568 434898 475610 435134
rect 475846 434898 475888 435134
rect 475568 434866 475888 434898
rect 506288 435454 506608 435486
rect 506288 435218 506330 435454
rect 506566 435218 506608 435454
rect 506288 435134 506608 435218
rect 506288 434898 506330 435134
rect 506566 434898 506608 435134
rect 506288 434866 506608 434898
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 91568 403954 91888 403986
rect 91568 403718 91610 403954
rect 91846 403718 91888 403954
rect 91568 403634 91888 403718
rect 91568 403398 91610 403634
rect 91846 403398 91888 403634
rect 91568 403366 91888 403398
rect 122288 403954 122608 403986
rect 122288 403718 122330 403954
rect 122566 403718 122608 403954
rect 122288 403634 122608 403718
rect 122288 403398 122330 403634
rect 122566 403398 122608 403634
rect 122288 403366 122608 403398
rect 153008 403954 153328 403986
rect 153008 403718 153050 403954
rect 153286 403718 153328 403954
rect 153008 403634 153328 403718
rect 153008 403398 153050 403634
rect 153286 403398 153328 403634
rect 153008 403366 153328 403398
rect 183728 403954 184048 403986
rect 183728 403718 183770 403954
rect 184006 403718 184048 403954
rect 183728 403634 184048 403718
rect 183728 403398 183770 403634
rect 184006 403398 184048 403634
rect 183728 403366 184048 403398
rect 214448 403954 214768 403986
rect 214448 403718 214490 403954
rect 214726 403718 214768 403954
rect 214448 403634 214768 403718
rect 214448 403398 214490 403634
rect 214726 403398 214768 403634
rect 214448 403366 214768 403398
rect 245168 403954 245488 403986
rect 245168 403718 245210 403954
rect 245446 403718 245488 403954
rect 245168 403634 245488 403718
rect 245168 403398 245210 403634
rect 245446 403398 245488 403634
rect 245168 403366 245488 403398
rect 275888 403954 276208 403986
rect 275888 403718 275930 403954
rect 276166 403718 276208 403954
rect 275888 403634 276208 403718
rect 275888 403398 275930 403634
rect 276166 403398 276208 403634
rect 275888 403366 276208 403398
rect 306608 403954 306928 403986
rect 306608 403718 306650 403954
rect 306886 403718 306928 403954
rect 306608 403634 306928 403718
rect 306608 403398 306650 403634
rect 306886 403398 306928 403634
rect 306608 403366 306928 403398
rect 337328 403954 337648 403986
rect 337328 403718 337370 403954
rect 337606 403718 337648 403954
rect 337328 403634 337648 403718
rect 337328 403398 337370 403634
rect 337606 403398 337648 403634
rect 337328 403366 337648 403398
rect 368048 403954 368368 403986
rect 368048 403718 368090 403954
rect 368326 403718 368368 403954
rect 368048 403634 368368 403718
rect 368048 403398 368090 403634
rect 368326 403398 368368 403634
rect 368048 403366 368368 403398
rect 398768 403954 399088 403986
rect 398768 403718 398810 403954
rect 399046 403718 399088 403954
rect 398768 403634 399088 403718
rect 398768 403398 398810 403634
rect 399046 403398 399088 403634
rect 398768 403366 399088 403398
rect 429488 403954 429808 403986
rect 429488 403718 429530 403954
rect 429766 403718 429808 403954
rect 429488 403634 429808 403718
rect 429488 403398 429530 403634
rect 429766 403398 429808 403634
rect 429488 403366 429808 403398
rect 460208 403954 460528 403986
rect 460208 403718 460250 403954
rect 460486 403718 460528 403954
rect 460208 403634 460528 403718
rect 460208 403398 460250 403634
rect 460486 403398 460528 403634
rect 460208 403366 460528 403398
rect 490928 403954 491248 403986
rect 490928 403718 490970 403954
rect 491206 403718 491248 403954
rect 490928 403634 491248 403718
rect 490928 403398 490970 403634
rect 491206 403398 491248 403634
rect 490928 403366 491248 403398
rect 76208 399454 76528 399486
rect 76208 399218 76250 399454
rect 76486 399218 76528 399454
rect 76208 399134 76528 399218
rect 76208 398898 76250 399134
rect 76486 398898 76528 399134
rect 76208 398866 76528 398898
rect 106928 399454 107248 399486
rect 106928 399218 106970 399454
rect 107206 399218 107248 399454
rect 106928 399134 107248 399218
rect 106928 398898 106970 399134
rect 107206 398898 107248 399134
rect 106928 398866 107248 398898
rect 137648 399454 137968 399486
rect 137648 399218 137690 399454
rect 137926 399218 137968 399454
rect 137648 399134 137968 399218
rect 137648 398898 137690 399134
rect 137926 398898 137968 399134
rect 137648 398866 137968 398898
rect 168368 399454 168688 399486
rect 168368 399218 168410 399454
rect 168646 399218 168688 399454
rect 168368 399134 168688 399218
rect 168368 398898 168410 399134
rect 168646 398898 168688 399134
rect 168368 398866 168688 398898
rect 199088 399454 199408 399486
rect 199088 399218 199130 399454
rect 199366 399218 199408 399454
rect 199088 399134 199408 399218
rect 199088 398898 199130 399134
rect 199366 398898 199408 399134
rect 199088 398866 199408 398898
rect 229808 399454 230128 399486
rect 229808 399218 229850 399454
rect 230086 399218 230128 399454
rect 229808 399134 230128 399218
rect 229808 398898 229850 399134
rect 230086 398898 230128 399134
rect 229808 398866 230128 398898
rect 260528 399454 260848 399486
rect 260528 399218 260570 399454
rect 260806 399218 260848 399454
rect 260528 399134 260848 399218
rect 260528 398898 260570 399134
rect 260806 398898 260848 399134
rect 260528 398866 260848 398898
rect 291248 399454 291568 399486
rect 291248 399218 291290 399454
rect 291526 399218 291568 399454
rect 291248 399134 291568 399218
rect 291248 398898 291290 399134
rect 291526 398898 291568 399134
rect 291248 398866 291568 398898
rect 321968 399454 322288 399486
rect 321968 399218 322010 399454
rect 322246 399218 322288 399454
rect 321968 399134 322288 399218
rect 321968 398898 322010 399134
rect 322246 398898 322288 399134
rect 321968 398866 322288 398898
rect 352688 399454 353008 399486
rect 352688 399218 352730 399454
rect 352966 399218 353008 399454
rect 352688 399134 353008 399218
rect 352688 398898 352730 399134
rect 352966 398898 353008 399134
rect 352688 398866 353008 398898
rect 383408 399454 383728 399486
rect 383408 399218 383450 399454
rect 383686 399218 383728 399454
rect 383408 399134 383728 399218
rect 383408 398898 383450 399134
rect 383686 398898 383728 399134
rect 383408 398866 383728 398898
rect 414128 399454 414448 399486
rect 414128 399218 414170 399454
rect 414406 399218 414448 399454
rect 414128 399134 414448 399218
rect 414128 398898 414170 399134
rect 414406 398898 414448 399134
rect 414128 398866 414448 398898
rect 444848 399454 445168 399486
rect 444848 399218 444890 399454
rect 445126 399218 445168 399454
rect 444848 399134 445168 399218
rect 444848 398898 444890 399134
rect 445126 398898 445168 399134
rect 444848 398866 445168 398898
rect 475568 399454 475888 399486
rect 475568 399218 475610 399454
rect 475846 399218 475888 399454
rect 475568 399134 475888 399218
rect 475568 398898 475610 399134
rect 475846 398898 475888 399134
rect 475568 398866 475888 398898
rect 506288 399454 506608 399486
rect 506288 399218 506330 399454
rect 506566 399218 506608 399454
rect 506288 399134 506608 399218
rect 506288 398898 506330 399134
rect 506566 398898 506608 399134
rect 506288 398866 506608 398898
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 91568 367954 91888 367986
rect 91568 367718 91610 367954
rect 91846 367718 91888 367954
rect 91568 367634 91888 367718
rect 91568 367398 91610 367634
rect 91846 367398 91888 367634
rect 91568 367366 91888 367398
rect 122288 367954 122608 367986
rect 122288 367718 122330 367954
rect 122566 367718 122608 367954
rect 122288 367634 122608 367718
rect 122288 367398 122330 367634
rect 122566 367398 122608 367634
rect 122288 367366 122608 367398
rect 153008 367954 153328 367986
rect 153008 367718 153050 367954
rect 153286 367718 153328 367954
rect 153008 367634 153328 367718
rect 153008 367398 153050 367634
rect 153286 367398 153328 367634
rect 153008 367366 153328 367398
rect 183728 367954 184048 367986
rect 183728 367718 183770 367954
rect 184006 367718 184048 367954
rect 183728 367634 184048 367718
rect 183728 367398 183770 367634
rect 184006 367398 184048 367634
rect 183728 367366 184048 367398
rect 214448 367954 214768 367986
rect 214448 367718 214490 367954
rect 214726 367718 214768 367954
rect 214448 367634 214768 367718
rect 214448 367398 214490 367634
rect 214726 367398 214768 367634
rect 214448 367366 214768 367398
rect 245168 367954 245488 367986
rect 245168 367718 245210 367954
rect 245446 367718 245488 367954
rect 245168 367634 245488 367718
rect 245168 367398 245210 367634
rect 245446 367398 245488 367634
rect 245168 367366 245488 367398
rect 275888 367954 276208 367986
rect 275888 367718 275930 367954
rect 276166 367718 276208 367954
rect 275888 367634 276208 367718
rect 275888 367398 275930 367634
rect 276166 367398 276208 367634
rect 275888 367366 276208 367398
rect 306608 367954 306928 367986
rect 306608 367718 306650 367954
rect 306886 367718 306928 367954
rect 306608 367634 306928 367718
rect 306608 367398 306650 367634
rect 306886 367398 306928 367634
rect 306608 367366 306928 367398
rect 337328 367954 337648 367986
rect 337328 367718 337370 367954
rect 337606 367718 337648 367954
rect 337328 367634 337648 367718
rect 337328 367398 337370 367634
rect 337606 367398 337648 367634
rect 337328 367366 337648 367398
rect 368048 367954 368368 367986
rect 368048 367718 368090 367954
rect 368326 367718 368368 367954
rect 368048 367634 368368 367718
rect 368048 367398 368090 367634
rect 368326 367398 368368 367634
rect 368048 367366 368368 367398
rect 398768 367954 399088 367986
rect 398768 367718 398810 367954
rect 399046 367718 399088 367954
rect 398768 367634 399088 367718
rect 398768 367398 398810 367634
rect 399046 367398 399088 367634
rect 398768 367366 399088 367398
rect 429488 367954 429808 367986
rect 429488 367718 429530 367954
rect 429766 367718 429808 367954
rect 429488 367634 429808 367718
rect 429488 367398 429530 367634
rect 429766 367398 429808 367634
rect 429488 367366 429808 367398
rect 460208 367954 460528 367986
rect 460208 367718 460250 367954
rect 460486 367718 460528 367954
rect 460208 367634 460528 367718
rect 460208 367398 460250 367634
rect 460486 367398 460528 367634
rect 460208 367366 460528 367398
rect 490928 367954 491248 367986
rect 490928 367718 490970 367954
rect 491206 367718 491248 367954
rect 490928 367634 491248 367718
rect 490928 367398 490970 367634
rect 491206 367398 491248 367634
rect 490928 367366 491248 367398
rect 76208 363454 76528 363486
rect 76208 363218 76250 363454
rect 76486 363218 76528 363454
rect 76208 363134 76528 363218
rect 76208 362898 76250 363134
rect 76486 362898 76528 363134
rect 76208 362866 76528 362898
rect 106928 363454 107248 363486
rect 106928 363218 106970 363454
rect 107206 363218 107248 363454
rect 106928 363134 107248 363218
rect 106928 362898 106970 363134
rect 107206 362898 107248 363134
rect 106928 362866 107248 362898
rect 137648 363454 137968 363486
rect 137648 363218 137690 363454
rect 137926 363218 137968 363454
rect 137648 363134 137968 363218
rect 137648 362898 137690 363134
rect 137926 362898 137968 363134
rect 137648 362866 137968 362898
rect 168368 363454 168688 363486
rect 168368 363218 168410 363454
rect 168646 363218 168688 363454
rect 168368 363134 168688 363218
rect 168368 362898 168410 363134
rect 168646 362898 168688 363134
rect 168368 362866 168688 362898
rect 199088 363454 199408 363486
rect 199088 363218 199130 363454
rect 199366 363218 199408 363454
rect 199088 363134 199408 363218
rect 199088 362898 199130 363134
rect 199366 362898 199408 363134
rect 199088 362866 199408 362898
rect 229808 363454 230128 363486
rect 229808 363218 229850 363454
rect 230086 363218 230128 363454
rect 229808 363134 230128 363218
rect 229808 362898 229850 363134
rect 230086 362898 230128 363134
rect 229808 362866 230128 362898
rect 260528 363454 260848 363486
rect 260528 363218 260570 363454
rect 260806 363218 260848 363454
rect 260528 363134 260848 363218
rect 260528 362898 260570 363134
rect 260806 362898 260848 363134
rect 260528 362866 260848 362898
rect 291248 363454 291568 363486
rect 291248 363218 291290 363454
rect 291526 363218 291568 363454
rect 291248 363134 291568 363218
rect 291248 362898 291290 363134
rect 291526 362898 291568 363134
rect 291248 362866 291568 362898
rect 321968 363454 322288 363486
rect 321968 363218 322010 363454
rect 322246 363218 322288 363454
rect 321968 363134 322288 363218
rect 321968 362898 322010 363134
rect 322246 362898 322288 363134
rect 321968 362866 322288 362898
rect 352688 363454 353008 363486
rect 352688 363218 352730 363454
rect 352966 363218 353008 363454
rect 352688 363134 353008 363218
rect 352688 362898 352730 363134
rect 352966 362898 353008 363134
rect 352688 362866 353008 362898
rect 383408 363454 383728 363486
rect 383408 363218 383450 363454
rect 383686 363218 383728 363454
rect 383408 363134 383728 363218
rect 383408 362898 383450 363134
rect 383686 362898 383728 363134
rect 383408 362866 383728 362898
rect 414128 363454 414448 363486
rect 414128 363218 414170 363454
rect 414406 363218 414448 363454
rect 414128 363134 414448 363218
rect 414128 362898 414170 363134
rect 414406 362898 414448 363134
rect 414128 362866 414448 362898
rect 444848 363454 445168 363486
rect 444848 363218 444890 363454
rect 445126 363218 445168 363454
rect 444848 363134 445168 363218
rect 444848 362898 444890 363134
rect 445126 362898 445168 363134
rect 444848 362866 445168 362898
rect 475568 363454 475888 363486
rect 475568 363218 475610 363454
rect 475846 363218 475888 363454
rect 475568 363134 475888 363218
rect 475568 362898 475610 363134
rect 475846 362898 475888 363134
rect 475568 362866 475888 362898
rect 506288 363454 506608 363486
rect 506288 363218 506330 363454
rect 506566 363218 506608 363454
rect 506288 363134 506608 363218
rect 506288 362898 506330 363134
rect 506566 362898 506608 363134
rect 506288 362866 506608 362898
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 91568 331954 91888 331986
rect 91568 331718 91610 331954
rect 91846 331718 91888 331954
rect 91568 331634 91888 331718
rect 91568 331398 91610 331634
rect 91846 331398 91888 331634
rect 91568 331366 91888 331398
rect 122288 331954 122608 331986
rect 122288 331718 122330 331954
rect 122566 331718 122608 331954
rect 122288 331634 122608 331718
rect 122288 331398 122330 331634
rect 122566 331398 122608 331634
rect 122288 331366 122608 331398
rect 153008 331954 153328 331986
rect 153008 331718 153050 331954
rect 153286 331718 153328 331954
rect 153008 331634 153328 331718
rect 153008 331398 153050 331634
rect 153286 331398 153328 331634
rect 153008 331366 153328 331398
rect 183728 331954 184048 331986
rect 183728 331718 183770 331954
rect 184006 331718 184048 331954
rect 183728 331634 184048 331718
rect 183728 331398 183770 331634
rect 184006 331398 184048 331634
rect 183728 331366 184048 331398
rect 214448 331954 214768 331986
rect 214448 331718 214490 331954
rect 214726 331718 214768 331954
rect 214448 331634 214768 331718
rect 214448 331398 214490 331634
rect 214726 331398 214768 331634
rect 214448 331366 214768 331398
rect 245168 331954 245488 331986
rect 245168 331718 245210 331954
rect 245446 331718 245488 331954
rect 245168 331634 245488 331718
rect 245168 331398 245210 331634
rect 245446 331398 245488 331634
rect 245168 331366 245488 331398
rect 275888 331954 276208 331986
rect 275888 331718 275930 331954
rect 276166 331718 276208 331954
rect 275888 331634 276208 331718
rect 275888 331398 275930 331634
rect 276166 331398 276208 331634
rect 275888 331366 276208 331398
rect 306608 331954 306928 331986
rect 306608 331718 306650 331954
rect 306886 331718 306928 331954
rect 306608 331634 306928 331718
rect 306608 331398 306650 331634
rect 306886 331398 306928 331634
rect 306608 331366 306928 331398
rect 337328 331954 337648 331986
rect 337328 331718 337370 331954
rect 337606 331718 337648 331954
rect 337328 331634 337648 331718
rect 337328 331398 337370 331634
rect 337606 331398 337648 331634
rect 337328 331366 337648 331398
rect 368048 331954 368368 331986
rect 368048 331718 368090 331954
rect 368326 331718 368368 331954
rect 368048 331634 368368 331718
rect 368048 331398 368090 331634
rect 368326 331398 368368 331634
rect 368048 331366 368368 331398
rect 398768 331954 399088 331986
rect 398768 331718 398810 331954
rect 399046 331718 399088 331954
rect 398768 331634 399088 331718
rect 398768 331398 398810 331634
rect 399046 331398 399088 331634
rect 398768 331366 399088 331398
rect 429488 331954 429808 331986
rect 429488 331718 429530 331954
rect 429766 331718 429808 331954
rect 429488 331634 429808 331718
rect 429488 331398 429530 331634
rect 429766 331398 429808 331634
rect 429488 331366 429808 331398
rect 460208 331954 460528 331986
rect 460208 331718 460250 331954
rect 460486 331718 460528 331954
rect 460208 331634 460528 331718
rect 460208 331398 460250 331634
rect 460486 331398 460528 331634
rect 460208 331366 460528 331398
rect 490928 331954 491248 331986
rect 490928 331718 490970 331954
rect 491206 331718 491248 331954
rect 490928 331634 491248 331718
rect 490928 331398 490970 331634
rect 491206 331398 491248 331634
rect 490928 331366 491248 331398
rect 76208 327454 76528 327486
rect 76208 327218 76250 327454
rect 76486 327218 76528 327454
rect 76208 327134 76528 327218
rect 76208 326898 76250 327134
rect 76486 326898 76528 327134
rect 76208 326866 76528 326898
rect 106928 327454 107248 327486
rect 106928 327218 106970 327454
rect 107206 327218 107248 327454
rect 106928 327134 107248 327218
rect 106928 326898 106970 327134
rect 107206 326898 107248 327134
rect 106928 326866 107248 326898
rect 137648 327454 137968 327486
rect 137648 327218 137690 327454
rect 137926 327218 137968 327454
rect 137648 327134 137968 327218
rect 137648 326898 137690 327134
rect 137926 326898 137968 327134
rect 137648 326866 137968 326898
rect 168368 327454 168688 327486
rect 168368 327218 168410 327454
rect 168646 327218 168688 327454
rect 168368 327134 168688 327218
rect 168368 326898 168410 327134
rect 168646 326898 168688 327134
rect 168368 326866 168688 326898
rect 199088 327454 199408 327486
rect 199088 327218 199130 327454
rect 199366 327218 199408 327454
rect 199088 327134 199408 327218
rect 199088 326898 199130 327134
rect 199366 326898 199408 327134
rect 199088 326866 199408 326898
rect 229808 327454 230128 327486
rect 229808 327218 229850 327454
rect 230086 327218 230128 327454
rect 229808 327134 230128 327218
rect 229808 326898 229850 327134
rect 230086 326898 230128 327134
rect 229808 326866 230128 326898
rect 260528 327454 260848 327486
rect 260528 327218 260570 327454
rect 260806 327218 260848 327454
rect 260528 327134 260848 327218
rect 260528 326898 260570 327134
rect 260806 326898 260848 327134
rect 260528 326866 260848 326898
rect 291248 327454 291568 327486
rect 291248 327218 291290 327454
rect 291526 327218 291568 327454
rect 291248 327134 291568 327218
rect 291248 326898 291290 327134
rect 291526 326898 291568 327134
rect 291248 326866 291568 326898
rect 321968 327454 322288 327486
rect 321968 327218 322010 327454
rect 322246 327218 322288 327454
rect 321968 327134 322288 327218
rect 321968 326898 322010 327134
rect 322246 326898 322288 327134
rect 321968 326866 322288 326898
rect 352688 327454 353008 327486
rect 352688 327218 352730 327454
rect 352966 327218 353008 327454
rect 352688 327134 353008 327218
rect 352688 326898 352730 327134
rect 352966 326898 353008 327134
rect 352688 326866 353008 326898
rect 383408 327454 383728 327486
rect 383408 327218 383450 327454
rect 383686 327218 383728 327454
rect 383408 327134 383728 327218
rect 383408 326898 383450 327134
rect 383686 326898 383728 327134
rect 383408 326866 383728 326898
rect 414128 327454 414448 327486
rect 414128 327218 414170 327454
rect 414406 327218 414448 327454
rect 414128 327134 414448 327218
rect 414128 326898 414170 327134
rect 414406 326898 414448 327134
rect 414128 326866 414448 326898
rect 444848 327454 445168 327486
rect 444848 327218 444890 327454
rect 445126 327218 445168 327454
rect 444848 327134 445168 327218
rect 444848 326898 444890 327134
rect 445126 326898 445168 327134
rect 444848 326866 445168 326898
rect 475568 327454 475888 327486
rect 475568 327218 475610 327454
rect 475846 327218 475888 327454
rect 475568 327134 475888 327218
rect 475568 326898 475610 327134
rect 475846 326898 475888 327134
rect 475568 326866 475888 326898
rect 506288 327454 506608 327486
rect 506288 327218 506330 327454
rect 506566 327218 506608 327454
rect 506288 327134 506608 327218
rect 506288 326898 506330 327134
rect 506566 326898 506608 327134
rect 506288 326866 506608 326898
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 91568 295954 91888 295986
rect 91568 295718 91610 295954
rect 91846 295718 91888 295954
rect 91568 295634 91888 295718
rect 91568 295398 91610 295634
rect 91846 295398 91888 295634
rect 91568 295366 91888 295398
rect 122288 295954 122608 295986
rect 122288 295718 122330 295954
rect 122566 295718 122608 295954
rect 122288 295634 122608 295718
rect 122288 295398 122330 295634
rect 122566 295398 122608 295634
rect 122288 295366 122608 295398
rect 153008 295954 153328 295986
rect 153008 295718 153050 295954
rect 153286 295718 153328 295954
rect 153008 295634 153328 295718
rect 153008 295398 153050 295634
rect 153286 295398 153328 295634
rect 153008 295366 153328 295398
rect 183728 295954 184048 295986
rect 183728 295718 183770 295954
rect 184006 295718 184048 295954
rect 183728 295634 184048 295718
rect 183728 295398 183770 295634
rect 184006 295398 184048 295634
rect 183728 295366 184048 295398
rect 214448 295954 214768 295986
rect 214448 295718 214490 295954
rect 214726 295718 214768 295954
rect 214448 295634 214768 295718
rect 214448 295398 214490 295634
rect 214726 295398 214768 295634
rect 214448 295366 214768 295398
rect 245168 295954 245488 295986
rect 245168 295718 245210 295954
rect 245446 295718 245488 295954
rect 245168 295634 245488 295718
rect 245168 295398 245210 295634
rect 245446 295398 245488 295634
rect 245168 295366 245488 295398
rect 275888 295954 276208 295986
rect 275888 295718 275930 295954
rect 276166 295718 276208 295954
rect 275888 295634 276208 295718
rect 275888 295398 275930 295634
rect 276166 295398 276208 295634
rect 275888 295366 276208 295398
rect 306608 295954 306928 295986
rect 306608 295718 306650 295954
rect 306886 295718 306928 295954
rect 306608 295634 306928 295718
rect 306608 295398 306650 295634
rect 306886 295398 306928 295634
rect 306608 295366 306928 295398
rect 337328 295954 337648 295986
rect 337328 295718 337370 295954
rect 337606 295718 337648 295954
rect 337328 295634 337648 295718
rect 337328 295398 337370 295634
rect 337606 295398 337648 295634
rect 337328 295366 337648 295398
rect 368048 295954 368368 295986
rect 368048 295718 368090 295954
rect 368326 295718 368368 295954
rect 368048 295634 368368 295718
rect 368048 295398 368090 295634
rect 368326 295398 368368 295634
rect 368048 295366 368368 295398
rect 398768 295954 399088 295986
rect 398768 295718 398810 295954
rect 399046 295718 399088 295954
rect 398768 295634 399088 295718
rect 398768 295398 398810 295634
rect 399046 295398 399088 295634
rect 398768 295366 399088 295398
rect 429488 295954 429808 295986
rect 429488 295718 429530 295954
rect 429766 295718 429808 295954
rect 429488 295634 429808 295718
rect 429488 295398 429530 295634
rect 429766 295398 429808 295634
rect 429488 295366 429808 295398
rect 460208 295954 460528 295986
rect 460208 295718 460250 295954
rect 460486 295718 460528 295954
rect 460208 295634 460528 295718
rect 460208 295398 460250 295634
rect 460486 295398 460528 295634
rect 460208 295366 460528 295398
rect 490928 295954 491248 295986
rect 490928 295718 490970 295954
rect 491206 295718 491248 295954
rect 490928 295634 491248 295718
rect 490928 295398 490970 295634
rect 491206 295398 491248 295634
rect 490928 295366 491248 295398
rect 76208 291454 76528 291486
rect 76208 291218 76250 291454
rect 76486 291218 76528 291454
rect 76208 291134 76528 291218
rect 76208 290898 76250 291134
rect 76486 290898 76528 291134
rect 76208 290866 76528 290898
rect 106928 291454 107248 291486
rect 106928 291218 106970 291454
rect 107206 291218 107248 291454
rect 106928 291134 107248 291218
rect 106928 290898 106970 291134
rect 107206 290898 107248 291134
rect 106928 290866 107248 290898
rect 137648 291454 137968 291486
rect 137648 291218 137690 291454
rect 137926 291218 137968 291454
rect 137648 291134 137968 291218
rect 137648 290898 137690 291134
rect 137926 290898 137968 291134
rect 137648 290866 137968 290898
rect 168368 291454 168688 291486
rect 168368 291218 168410 291454
rect 168646 291218 168688 291454
rect 168368 291134 168688 291218
rect 168368 290898 168410 291134
rect 168646 290898 168688 291134
rect 168368 290866 168688 290898
rect 199088 291454 199408 291486
rect 199088 291218 199130 291454
rect 199366 291218 199408 291454
rect 199088 291134 199408 291218
rect 199088 290898 199130 291134
rect 199366 290898 199408 291134
rect 199088 290866 199408 290898
rect 229808 291454 230128 291486
rect 229808 291218 229850 291454
rect 230086 291218 230128 291454
rect 229808 291134 230128 291218
rect 229808 290898 229850 291134
rect 230086 290898 230128 291134
rect 229808 290866 230128 290898
rect 260528 291454 260848 291486
rect 260528 291218 260570 291454
rect 260806 291218 260848 291454
rect 260528 291134 260848 291218
rect 260528 290898 260570 291134
rect 260806 290898 260848 291134
rect 260528 290866 260848 290898
rect 291248 291454 291568 291486
rect 291248 291218 291290 291454
rect 291526 291218 291568 291454
rect 291248 291134 291568 291218
rect 291248 290898 291290 291134
rect 291526 290898 291568 291134
rect 291248 290866 291568 290898
rect 321968 291454 322288 291486
rect 321968 291218 322010 291454
rect 322246 291218 322288 291454
rect 321968 291134 322288 291218
rect 321968 290898 322010 291134
rect 322246 290898 322288 291134
rect 321968 290866 322288 290898
rect 352688 291454 353008 291486
rect 352688 291218 352730 291454
rect 352966 291218 353008 291454
rect 352688 291134 353008 291218
rect 352688 290898 352730 291134
rect 352966 290898 353008 291134
rect 352688 290866 353008 290898
rect 383408 291454 383728 291486
rect 383408 291218 383450 291454
rect 383686 291218 383728 291454
rect 383408 291134 383728 291218
rect 383408 290898 383450 291134
rect 383686 290898 383728 291134
rect 383408 290866 383728 290898
rect 414128 291454 414448 291486
rect 414128 291218 414170 291454
rect 414406 291218 414448 291454
rect 414128 291134 414448 291218
rect 414128 290898 414170 291134
rect 414406 290898 414448 291134
rect 414128 290866 414448 290898
rect 444848 291454 445168 291486
rect 444848 291218 444890 291454
rect 445126 291218 445168 291454
rect 444848 291134 445168 291218
rect 444848 290898 444890 291134
rect 445126 290898 445168 291134
rect 444848 290866 445168 290898
rect 475568 291454 475888 291486
rect 475568 291218 475610 291454
rect 475846 291218 475888 291454
rect 475568 291134 475888 291218
rect 475568 290898 475610 291134
rect 475846 290898 475888 291134
rect 475568 290866 475888 290898
rect 506288 291454 506608 291486
rect 506288 291218 506330 291454
rect 506566 291218 506608 291454
rect 506288 291134 506608 291218
rect 506288 290898 506330 291134
rect 506566 290898 506608 291134
rect 506288 290866 506608 290898
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 91568 259954 91888 259986
rect 91568 259718 91610 259954
rect 91846 259718 91888 259954
rect 91568 259634 91888 259718
rect 91568 259398 91610 259634
rect 91846 259398 91888 259634
rect 91568 259366 91888 259398
rect 122288 259954 122608 259986
rect 122288 259718 122330 259954
rect 122566 259718 122608 259954
rect 122288 259634 122608 259718
rect 122288 259398 122330 259634
rect 122566 259398 122608 259634
rect 122288 259366 122608 259398
rect 153008 259954 153328 259986
rect 153008 259718 153050 259954
rect 153286 259718 153328 259954
rect 153008 259634 153328 259718
rect 153008 259398 153050 259634
rect 153286 259398 153328 259634
rect 153008 259366 153328 259398
rect 183728 259954 184048 259986
rect 183728 259718 183770 259954
rect 184006 259718 184048 259954
rect 183728 259634 184048 259718
rect 183728 259398 183770 259634
rect 184006 259398 184048 259634
rect 183728 259366 184048 259398
rect 214448 259954 214768 259986
rect 214448 259718 214490 259954
rect 214726 259718 214768 259954
rect 214448 259634 214768 259718
rect 214448 259398 214490 259634
rect 214726 259398 214768 259634
rect 214448 259366 214768 259398
rect 245168 259954 245488 259986
rect 245168 259718 245210 259954
rect 245446 259718 245488 259954
rect 245168 259634 245488 259718
rect 245168 259398 245210 259634
rect 245446 259398 245488 259634
rect 245168 259366 245488 259398
rect 275888 259954 276208 259986
rect 275888 259718 275930 259954
rect 276166 259718 276208 259954
rect 275888 259634 276208 259718
rect 275888 259398 275930 259634
rect 276166 259398 276208 259634
rect 275888 259366 276208 259398
rect 306608 259954 306928 259986
rect 306608 259718 306650 259954
rect 306886 259718 306928 259954
rect 306608 259634 306928 259718
rect 306608 259398 306650 259634
rect 306886 259398 306928 259634
rect 306608 259366 306928 259398
rect 337328 259954 337648 259986
rect 337328 259718 337370 259954
rect 337606 259718 337648 259954
rect 337328 259634 337648 259718
rect 337328 259398 337370 259634
rect 337606 259398 337648 259634
rect 337328 259366 337648 259398
rect 368048 259954 368368 259986
rect 368048 259718 368090 259954
rect 368326 259718 368368 259954
rect 368048 259634 368368 259718
rect 368048 259398 368090 259634
rect 368326 259398 368368 259634
rect 368048 259366 368368 259398
rect 398768 259954 399088 259986
rect 398768 259718 398810 259954
rect 399046 259718 399088 259954
rect 398768 259634 399088 259718
rect 398768 259398 398810 259634
rect 399046 259398 399088 259634
rect 398768 259366 399088 259398
rect 429488 259954 429808 259986
rect 429488 259718 429530 259954
rect 429766 259718 429808 259954
rect 429488 259634 429808 259718
rect 429488 259398 429530 259634
rect 429766 259398 429808 259634
rect 429488 259366 429808 259398
rect 460208 259954 460528 259986
rect 460208 259718 460250 259954
rect 460486 259718 460528 259954
rect 460208 259634 460528 259718
rect 460208 259398 460250 259634
rect 460486 259398 460528 259634
rect 460208 259366 460528 259398
rect 490928 259954 491248 259986
rect 490928 259718 490970 259954
rect 491206 259718 491248 259954
rect 490928 259634 491248 259718
rect 490928 259398 490970 259634
rect 491206 259398 491248 259634
rect 490928 259366 491248 259398
rect 76208 255454 76528 255486
rect 76208 255218 76250 255454
rect 76486 255218 76528 255454
rect 76208 255134 76528 255218
rect 76208 254898 76250 255134
rect 76486 254898 76528 255134
rect 76208 254866 76528 254898
rect 106928 255454 107248 255486
rect 106928 255218 106970 255454
rect 107206 255218 107248 255454
rect 106928 255134 107248 255218
rect 106928 254898 106970 255134
rect 107206 254898 107248 255134
rect 106928 254866 107248 254898
rect 137648 255454 137968 255486
rect 137648 255218 137690 255454
rect 137926 255218 137968 255454
rect 137648 255134 137968 255218
rect 137648 254898 137690 255134
rect 137926 254898 137968 255134
rect 137648 254866 137968 254898
rect 168368 255454 168688 255486
rect 168368 255218 168410 255454
rect 168646 255218 168688 255454
rect 168368 255134 168688 255218
rect 168368 254898 168410 255134
rect 168646 254898 168688 255134
rect 168368 254866 168688 254898
rect 199088 255454 199408 255486
rect 199088 255218 199130 255454
rect 199366 255218 199408 255454
rect 199088 255134 199408 255218
rect 199088 254898 199130 255134
rect 199366 254898 199408 255134
rect 199088 254866 199408 254898
rect 229808 255454 230128 255486
rect 229808 255218 229850 255454
rect 230086 255218 230128 255454
rect 229808 255134 230128 255218
rect 229808 254898 229850 255134
rect 230086 254898 230128 255134
rect 229808 254866 230128 254898
rect 260528 255454 260848 255486
rect 260528 255218 260570 255454
rect 260806 255218 260848 255454
rect 260528 255134 260848 255218
rect 260528 254898 260570 255134
rect 260806 254898 260848 255134
rect 260528 254866 260848 254898
rect 291248 255454 291568 255486
rect 291248 255218 291290 255454
rect 291526 255218 291568 255454
rect 291248 255134 291568 255218
rect 291248 254898 291290 255134
rect 291526 254898 291568 255134
rect 291248 254866 291568 254898
rect 321968 255454 322288 255486
rect 321968 255218 322010 255454
rect 322246 255218 322288 255454
rect 321968 255134 322288 255218
rect 321968 254898 322010 255134
rect 322246 254898 322288 255134
rect 321968 254866 322288 254898
rect 352688 255454 353008 255486
rect 352688 255218 352730 255454
rect 352966 255218 353008 255454
rect 352688 255134 353008 255218
rect 352688 254898 352730 255134
rect 352966 254898 353008 255134
rect 352688 254866 353008 254898
rect 383408 255454 383728 255486
rect 383408 255218 383450 255454
rect 383686 255218 383728 255454
rect 383408 255134 383728 255218
rect 383408 254898 383450 255134
rect 383686 254898 383728 255134
rect 383408 254866 383728 254898
rect 414128 255454 414448 255486
rect 414128 255218 414170 255454
rect 414406 255218 414448 255454
rect 414128 255134 414448 255218
rect 414128 254898 414170 255134
rect 414406 254898 414448 255134
rect 414128 254866 414448 254898
rect 444848 255454 445168 255486
rect 444848 255218 444890 255454
rect 445126 255218 445168 255454
rect 444848 255134 445168 255218
rect 444848 254898 444890 255134
rect 445126 254898 445168 255134
rect 444848 254866 445168 254898
rect 475568 255454 475888 255486
rect 475568 255218 475610 255454
rect 475846 255218 475888 255454
rect 475568 255134 475888 255218
rect 475568 254898 475610 255134
rect 475846 254898 475888 255134
rect 475568 254866 475888 254898
rect 506288 255454 506608 255486
rect 506288 255218 506330 255454
rect 506566 255218 506608 255454
rect 506288 255134 506608 255218
rect 506288 254898 506330 255134
rect 506566 254898 506608 255134
rect 506288 254866 506608 254898
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 91568 223954 91888 223986
rect 91568 223718 91610 223954
rect 91846 223718 91888 223954
rect 91568 223634 91888 223718
rect 91568 223398 91610 223634
rect 91846 223398 91888 223634
rect 91568 223366 91888 223398
rect 122288 223954 122608 223986
rect 122288 223718 122330 223954
rect 122566 223718 122608 223954
rect 122288 223634 122608 223718
rect 122288 223398 122330 223634
rect 122566 223398 122608 223634
rect 122288 223366 122608 223398
rect 153008 223954 153328 223986
rect 153008 223718 153050 223954
rect 153286 223718 153328 223954
rect 153008 223634 153328 223718
rect 153008 223398 153050 223634
rect 153286 223398 153328 223634
rect 153008 223366 153328 223398
rect 183728 223954 184048 223986
rect 183728 223718 183770 223954
rect 184006 223718 184048 223954
rect 183728 223634 184048 223718
rect 183728 223398 183770 223634
rect 184006 223398 184048 223634
rect 183728 223366 184048 223398
rect 214448 223954 214768 223986
rect 214448 223718 214490 223954
rect 214726 223718 214768 223954
rect 214448 223634 214768 223718
rect 214448 223398 214490 223634
rect 214726 223398 214768 223634
rect 214448 223366 214768 223398
rect 245168 223954 245488 223986
rect 245168 223718 245210 223954
rect 245446 223718 245488 223954
rect 245168 223634 245488 223718
rect 245168 223398 245210 223634
rect 245446 223398 245488 223634
rect 245168 223366 245488 223398
rect 275888 223954 276208 223986
rect 275888 223718 275930 223954
rect 276166 223718 276208 223954
rect 275888 223634 276208 223718
rect 275888 223398 275930 223634
rect 276166 223398 276208 223634
rect 275888 223366 276208 223398
rect 306608 223954 306928 223986
rect 306608 223718 306650 223954
rect 306886 223718 306928 223954
rect 306608 223634 306928 223718
rect 306608 223398 306650 223634
rect 306886 223398 306928 223634
rect 306608 223366 306928 223398
rect 337328 223954 337648 223986
rect 337328 223718 337370 223954
rect 337606 223718 337648 223954
rect 337328 223634 337648 223718
rect 337328 223398 337370 223634
rect 337606 223398 337648 223634
rect 337328 223366 337648 223398
rect 368048 223954 368368 223986
rect 368048 223718 368090 223954
rect 368326 223718 368368 223954
rect 368048 223634 368368 223718
rect 368048 223398 368090 223634
rect 368326 223398 368368 223634
rect 368048 223366 368368 223398
rect 398768 223954 399088 223986
rect 398768 223718 398810 223954
rect 399046 223718 399088 223954
rect 398768 223634 399088 223718
rect 398768 223398 398810 223634
rect 399046 223398 399088 223634
rect 398768 223366 399088 223398
rect 429488 223954 429808 223986
rect 429488 223718 429530 223954
rect 429766 223718 429808 223954
rect 429488 223634 429808 223718
rect 429488 223398 429530 223634
rect 429766 223398 429808 223634
rect 429488 223366 429808 223398
rect 460208 223954 460528 223986
rect 460208 223718 460250 223954
rect 460486 223718 460528 223954
rect 460208 223634 460528 223718
rect 460208 223398 460250 223634
rect 460486 223398 460528 223634
rect 460208 223366 460528 223398
rect 490928 223954 491248 223986
rect 490928 223718 490970 223954
rect 491206 223718 491248 223954
rect 490928 223634 491248 223718
rect 490928 223398 490970 223634
rect 491206 223398 491248 223634
rect 490928 223366 491248 223398
rect 76208 219454 76528 219486
rect 76208 219218 76250 219454
rect 76486 219218 76528 219454
rect 76208 219134 76528 219218
rect 76208 218898 76250 219134
rect 76486 218898 76528 219134
rect 76208 218866 76528 218898
rect 106928 219454 107248 219486
rect 106928 219218 106970 219454
rect 107206 219218 107248 219454
rect 106928 219134 107248 219218
rect 106928 218898 106970 219134
rect 107206 218898 107248 219134
rect 106928 218866 107248 218898
rect 137648 219454 137968 219486
rect 137648 219218 137690 219454
rect 137926 219218 137968 219454
rect 137648 219134 137968 219218
rect 137648 218898 137690 219134
rect 137926 218898 137968 219134
rect 137648 218866 137968 218898
rect 168368 219454 168688 219486
rect 168368 219218 168410 219454
rect 168646 219218 168688 219454
rect 168368 219134 168688 219218
rect 168368 218898 168410 219134
rect 168646 218898 168688 219134
rect 168368 218866 168688 218898
rect 199088 219454 199408 219486
rect 199088 219218 199130 219454
rect 199366 219218 199408 219454
rect 199088 219134 199408 219218
rect 199088 218898 199130 219134
rect 199366 218898 199408 219134
rect 199088 218866 199408 218898
rect 229808 219454 230128 219486
rect 229808 219218 229850 219454
rect 230086 219218 230128 219454
rect 229808 219134 230128 219218
rect 229808 218898 229850 219134
rect 230086 218898 230128 219134
rect 229808 218866 230128 218898
rect 260528 219454 260848 219486
rect 260528 219218 260570 219454
rect 260806 219218 260848 219454
rect 260528 219134 260848 219218
rect 260528 218898 260570 219134
rect 260806 218898 260848 219134
rect 260528 218866 260848 218898
rect 291248 219454 291568 219486
rect 291248 219218 291290 219454
rect 291526 219218 291568 219454
rect 291248 219134 291568 219218
rect 291248 218898 291290 219134
rect 291526 218898 291568 219134
rect 291248 218866 291568 218898
rect 321968 219454 322288 219486
rect 321968 219218 322010 219454
rect 322246 219218 322288 219454
rect 321968 219134 322288 219218
rect 321968 218898 322010 219134
rect 322246 218898 322288 219134
rect 321968 218866 322288 218898
rect 352688 219454 353008 219486
rect 352688 219218 352730 219454
rect 352966 219218 353008 219454
rect 352688 219134 353008 219218
rect 352688 218898 352730 219134
rect 352966 218898 353008 219134
rect 352688 218866 353008 218898
rect 383408 219454 383728 219486
rect 383408 219218 383450 219454
rect 383686 219218 383728 219454
rect 383408 219134 383728 219218
rect 383408 218898 383450 219134
rect 383686 218898 383728 219134
rect 383408 218866 383728 218898
rect 414128 219454 414448 219486
rect 414128 219218 414170 219454
rect 414406 219218 414448 219454
rect 414128 219134 414448 219218
rect 414128 218898 414170 219134
rect 414406 218898 414448 219134
rect 414128 218866 414448 218898
rect 444848 219454 445168 219486
rect 444848 219218 444890 219454
rect 445126 219218 445168 219454
rect 444848 219134 445168 219218
rect 444848 218898 444890 219134
rect 445126 218898 445168 219134
rect 444848 218866 445168 218898
rect 475568 219454 475888 219486
rect 475568 219218 475610 219454
rect 475846 219218 475888 219454
rect 475568 219134 475888 219218
rect 475568 218898 475610 219134
rect 475846 218898 475888 219134
rect 475568 218866 475888 218898
rect 506288 219454 506608 219486
rect 506288 219218 506330 219454
rect 506566 219218 506608 219454
rect 506288 219134 506608 219218
rect 506288 218898 506330 219134
rect 506566 218898 506608 219134
rect 506288 218866 506608 218898
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 91568 187954 91888 187986
rect 91568 187718 91610 187954
rect 91846 187718 91888 187954
rect 91568 187634 91888 187718
rect 91568 187398 91610 187634
rect 91846 187398 91888 187634
rect 91568 187366 91888 187398
rect 122288 187954 122608 187986
rect 122288 187718 122330 187954
rect 122566 187718 122608 187954
rect 122288 187634 122608 187718
rect 122288 187398 122330 187634
rect 122566 187398 122608 187634
rect 122288 187366 122608 187398
rect 153008 187954 153328 187986
rect 153008 187718 153050 187954
rect 153286 187718 153328 187954
rect 153008 187634 153328 187718
rect 153008 187398 153050 187634
rect 153286 187398 153328 187634
rect 153008 187366 153328 187398
rect 183728 187954 184048 187986
rect 183728 187718 183770 187954
rect 184006 187718 184048 187954
rect 183728 187634 184048 187718
rect 183728 187398 183770 187634
rect 184006 187398 184048 187634
rect 183728 187366 184048 187398
rect 214448 187954 214768 187986
rect 214448 187718 214490 187954
rect 214726 187718 214768 187954
rect 214448 187634 214768 187718
rect 214448 187398 214490 187634
rect 214726 187398 214768 187634
rect 214448 187366 214768 187398
rect 245168 187954 245488 187986
rect 245168 187718 245210 187954
rect 245446 187718 245488 187954
rect 245168 187634 245488 187718
rect 245168 187398 245210 187634
rect 245446 187398 245488 187634
rect 245168 187366 245488 187398
rect 275888 187954 276208 187986
rect 275888 187718 275930 187954
rect 276166 187718 276208 187954
rect 275888 187634 276208 187718
rect 275888 187398 275930 187634
rect 276166 187398 276208 187634
rect 275888 187366 276208 187398
rect 306608 187954 306928 187986
rect 306608 187718 306650 187954
rect 306886 187718 306928 187954
rect 306608 187634 306928 187718
rect 306608 187398 306650 187634
rect 306886 187398 306928 187634
rect 306608 187366 306928 187398
rect 337328 187954 337648 187986
rect 337328 187718 337370 187954
rect 337606 187718 337648 187954
rect 337328 187634 337648 187718
rect 337328 187398 337370 187634
rect 337606 187398 337648 187634
rect 337328 187366 337648 187398
rect 368048 187954 368368 187986
rect 368048 187718 368090 187954
rect 368326 187718 368368 187954
rect 368048 187634 368368 187718
rect 368048 187398 368090 187634
rect 368326 187398 368368 187634
rect 368048 187366 368368 187398
rect 398768 187954 399088 187986
rect 398768 187718 398810 187954
rect 399046 187718 399088 187954
rect 398768 187634 399088 187718
rect 398768 187398 398810 187634
rect 399046 187398 399088 187634
rect 398768 187366 399088 187398
rect 429488 187954 429808 187986
rect 429488 187718 429530 187954
rect 429766 187718 429808 187954
rect 429488 187634 429808 187718
rect 429488 187398 429530 187634
rect 429766 187398 429808 187634
rect 429488 187366 429808 187398
rect 460208 187954 460528 187986
rect 460208 187718 460250 187954
rect 460486 187718 460528 187954
rect 460208 187634 460528 187718
rect 460208 187398 460250 187634
rect 460486 187398 460528 187634
rect 460208 187366 460528 187398
rect 490928 187954 491248 187986
rect 490928 187718 490970 187954
rect 491206 187718 491248 187954
rect 490928 187634 491248 187718
rect 490928 187398 490970 187634
rect 491206 187398 491248 187634
rect 490928 187366 491248 187398
rect 76208 183454 76528 183486
rect 76208 183218 76250 183454
rect 76486 183218 76528 183454
rect 76208 183134 76528 183218
rect 76208 182898 76250 183134
rect 76486 182898 76528 183134
rect 76208 182866 76528 182898
rect 106928 183454 107248 183486
rect 106928 183218 106970 183454
rect 107206 183218 107248 183454
rect 106928 183134 107248 183218
rect 106928 182898 106970 183134
rect 107206 182898 107248 183134
rect 106928 182866 107248 182898
rect 137648 183454 137968 183486
rect 137648 183218 137690 183454
rect 137926 183218 137968 183454
rect 137648 183134 137968 183218
rect 137648 182898 137690 183134
rect 137926 182898 137968 183134
rect 137648 182866 137968 182898
rect 168368 183454 168688 183486
rect 168368 183218 168410 183454
rect 168646 183218 168688 183454
rect 168368 183134 168688 183218
rect 168368 182898 168410 183134
rect 168646 182898 168688 183134
rect 168368 182866 168688 182898
rect 199088 183454 199408 183486
rect 199088 183218 199130 183454
rect 199366 183218 199408 183454
rect 199088 183134 199408 183218
rect 199088 182898 199130 183134
rect 199366 182898 199408 183134
rect 199088 182866 199408 182898
rect 229808 183454 230128 183486
rect 229808 183218 229850 183454
rect 230086 183218 230128 183454
rect 229808 183134 230128 183218
rect 229808 182898 229850 183134
rect 230086 182898 230128 183134
rect 229808 182866 230128 182898
rect 260528 183454 260848 183486
rect 260528 183218 260570 183454
rect 260806 183218 260848 183454
rect 260528 183134 260848 183218
rect 260528 182898 260570 183134
rect 260806 182898 260848 183134
rect 260528 182866 260848 182898
rect 291248 183454 291568 183486
rect 291248 183218 291290 183454
rect 291526 183218 291568 183454
rect 291248 183134 291568 183218
rect 291248 182898 291290 183134
rect 291526 182898 291568 183134
rect 291248 182866 291568 182898
rect 321968 183454 322288 183486
rect 321968 183218 322010 183454
rect 322246 183218 322288 183454
rect 321968 183134 322288 183218
rect 321968 182898 322010 183134
rect 322246 182898 322288 183134
rect 321968 182866 322288 182898
rect 352688 183454 353008 183486
rect 352688 183218 352730 183454
rect 352966 183218 353008 183454
rect 352688 183134 353008 183218
rect 352688 182898 352730 183134
rect 352966 182898 353008 183134
rect 352688 182866 353008 182898
rect 383408 183454 383728 183486
rect 383408 183218 383450 183454
rect 383686 183218 383728 183454
rect 383408 183134 383728 183218
rect 383408 182898 383450 183134
rect 383686 182898 383728 183134
rect 383408 182866 383728 182898
rect 414128 183454 414448 183486
rect 414128 183218 414170 183454
rect 414406 183218 414448 183454
rect 414128 183134 414448 183218
rect 414128 182898 414170 183134
rect 414406 182898 414448 183134
rect 414128 182866 414448 182898
rect 444848 183454 445168 183486
rect 444848 183218 444890 183454
rect 445126 183218 445168 183454
rect 444848 183134 445168 183218
rect 444848 182898 444890 183134
rect 445126 182898 445168 183134
rect 444848 182866 445168 182898
rect 475568 183454 475888 183486
rect 475568 183218 475610 183454
rect 475846 183218 475888 183454
rect 475568 183134 475888 183218
rect 475568 182898 475610 183134
rect 475846 182898 475888 183134
rect 475568 182866 475888 182898
rect 506288 183454 506608 183486
rect 506288 183218 506330 183454
rect 506566 183218 506608 183454
rect 506288 183134 506608 183218
rect 506288 182898 506330 183134
rect 506566 182898 506608 183134
rect 506288 182866 506608 182898
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 91568 151954 91888 151986
rect 91568 151718 91610 151954
rect 91846 151718 91888 151954
rect 91568 151634 91888 151718
rect 91568 151398 91610 151634
rect 91846 151398 91888 151634
rect 91568 151366 91888 151398
rect 122288 151954 122608 151986
rect 122288 151718 122330 151954
rect 122566 151718 122608 151954
rect 122288 151634 122608 151718
rect 122288 151398 122330 151634
rect 122566 151398 122608 151634
rect 122288 151366 122608 151398
rect 153008 151954 153328 151986
rect 153008 151718 153050 151954
rect 153286 151718 153328 151954
rect 153008 151634 153328 151718
rect 153008 151398 153050 151634
rect 153286 151398 153328 151634
rect 153008 151366 153328 151398
rect 183728 151954 184048 151986
rect 183728 151718 183770 151954
rect 184006 151718 184048 151954
rect 183728 151634 184048 151718
rect 183728 151398 183770 151634
rect 184006 151398 184048 151634
rect 183728 151366 184048 151398
rect 214448 151954 214768 151986
rect 214448 151718 214490 151954
rect 214726 151718 214768 151954
rect 214448 151634 214768 151718
rect 214448 151398 214490 151634
rect 214726 151398 214768 151634
rect 214448 151366 214768 151398
rect 245168 151954 245488 151986
rect 245168 151718 245210 151954
rect 245446 151718 245488 151954
rect 245168 151634 245488 151718
rect 245168 151398 245210 151634
rect 245446 151398 245488 151634
rect 245168 151366 245488 151398
rect 275888 151954 276208 151986
rect 275888 151718 275930 151954
rect 276166 151718 276208 151954
rect 275888 151634 276208 151718
rect 275888 151398 275930 151634
rect 276166 151398 276208 151634
rect 275888 151366 276208 151398
rect 306608 151954 306928 151986
rect 306608 151718 306650 151954
rect 306886 151718 306928 151954
rect 306608 151634 306928 151718
rect 306608 151398 306650 151634
rect 306886 151398 306928 151634
rect 306608 151366 306928 151398
rect 337328 151954 337648 151986
rect 337328 151718 337370 151954
rect 337606 151718 337648 151954
rect 337328 151634 337648 151718
rect 337328 151398 337370 151634
rect 337606 151398 337648 151634
rect 337328 151366 337648 151398
rect 368048 151954 368368 151986
rect 368048 151718 368090 151954
rect 368326 151718 368368 151954
rect 368048 151634 368368 151718
rect 368048 151398 368090 151634
rect 368326 151398 368368 151634
rect 368048 151366 368368 151398
rect 398768 151954 399088 151986
rect 398768 151718 398810 151954
rect 399046 151718 399088 151954
rect 398768 151634 399088 151718
rect 398768 151398 398810 151634
rect 399046 151398 399088 151634
rect 398768 151366 399088 151398
rect 429488 151954 429808 151986
rect 429488 151718 429530 151954
rect 429766 151718 429808 151954
rect 429488 151634 429808 151718
rect 429488 151398 429530 151634
rect 429766 151398 429808 151634
rect 429488 151366 429808 151398
rect 460208 151954 460528 151986
rect 460208 151718 460250 151954
rect 460486 151718 460528 151954
rect 460208 151634 460528 151718
rect 460208 151398 460250 151634
rect 460486 151398 460528 151634
rect 460208 151366 460528 151398
rect 490928 151954 491248 151986
rect 490928 151718 490970 151954
rect 491206 151718 491248 151954
rect 490928 151634 491248 151718
rect 490928 151398 490970 151634
rect 491206 151398 491248 151634
rect 490928 151366 491248 151398
rect 76208 147454 76528 147486
rect 76208 147218 76250 147454
rect 76486 147218 76528 147454
rect 76208 147134 76528 147218
rect 76208 146898 76250 147134
rect 76486 146898 76528 147134
rect 76208 146866 76528 146898
rect 106928 147454 107248 147486
rect 106928 147218 106970 147454
rect 107206 147218 107248 147454
rect 106928 147134 107248 147218
rect 106928 146898 106970 147134
rect 107206 146898 107248 147134
rect 106928 146866 107248 146898
rect 137648 147454 137968 147486
rect 137648 147218 137690 147454
rect 137926 147218 137968 147454
rect 137648 147134 137968 147218
rect 137648 146898 137690 147134
rect 137926 146898 137968 147134
rect 137648 146866 137968 146898
rect 168368 147454 168688 147486
rect 168368 147218 168410 147454
rect 168646 147218 168688 147454
rect 168368 147134 168688 147218
rect 168368 146898 168410 147134
rect 168646 146898 168688 147134
rect 168368 146866 168688 146898
rect 199088 147454 199408 147486
rect 199088 147218 199130 147454
rect 199366 147218 199408 147454
rect 199088 147134 199408 147218
rect 199088 146898 199130 147134
rect 199366 146898 199408 147134
rect 199088 146866 199408 146898
rect 229808 147454 230128 147486
rect 229808 147218 229850 147454
rect 230086 147218 230128 147454
rect 229808 147134 230128 147218
rect 229808 146898 229850 147134
rect 230086 146898 230128 147134
rect 229808 146866 230128 146898
rect 260528 147454 260848 147486
rect 260528 147218 260570 147454
rect 260806 147218 260848 147454
rect 260528 147134 260848 147218
rect 260528 146898 260570 147134
rect 260806 146898 260848 147134
rect 260528 146866 260848 146898
rect 291248 147454 291568 147486
rect 291248 147218 291290 147454
rect 291526 147218 291568 147454
rect 291248 147134 291568 147218
rect 291248 146898 291290 147134
rect 291526 146898 291568 147134
rect 291248 146866 291568 146898
rect 321968 147454 322288 147486
rect 321968 147218 322010 147454
rect 322246 147218 322288 147454
rect 321968 147134 322288 147218
rect 321968 146898 322010 147134
rect 322246 146898 322288 147134
rect 321968 146866 322288 146898
rect 352688 147454 353008 147486
rect 352688 147218 352730 147454
rect 352966 147218 353008 147454
rect 352688 147134 353008 147218
rect 352688 146898 352730 147134
rect 352966 146898 353008 147134
rect 352688 146866 353008 146898
rect 383408 147454 383728 147486
rect 383408 147218 383450 147454
rect 383686 147218 383728 147454
rect 383408 147134 383728 147218
rect 383408 146898 383450 147134
rect 383686 146898 383728 147134
rect 383408 146866 383728 146898
rect 414128 147454 414448 147486
rect 414128 147218 414170 147454
rect 414406 147218 414448 147454
rect 414128 147134 414448 147218
rect 414128 146898 414170 147134
rect 414406 146898 414448 147134
rect 414128 146866 414448 146898
rect 444848 147454 445168 147486
rect 444848 147218 444890 147454
rect 445126 147218 445168 147454
rect 444848 147134 445168 147218
rect 444848 146898 444890 147134
rect 445126 146898 445168 147134
rect 444848 146866 445168 146898
rect 475568 147454 475888 147486
rect 475568 147218 475610 147454
rect 475846 147218 475888 147454
rect 475568 147134 475888 147218
rect 475568 146898 475610 147134
rect 475846 146898 475888 147134
rect 475568 146866 475888 146898
rect 506288 147454 506608 147486
rect 506288 147218 506330 147454
rect 506566 147218 506608 147454
rect 506288 147134 506608 147218
rect 506288 146898 506330 147134
rect 506566 146898 506608 147134
rect 506288 146866 506608 146898
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 91568 115954 91888 115986
rect 91568 115718 91610 115954
rect 91846 115718 91888 115954
rect 91568 115634 91888 115718
rect 91568 115398 91610 115634
rect 91846 115398 91888 115634
rect 91568 115366 91888 115398
rect 122288 115954 122608 115986
rect 122288 115718 122330 115954
rect 122566 115718 122608 115954
rect 122288 115634 122608 115718
rect 122288 115398 122330 115634
rect 122566 115398 122608 115634
rect 122288 115366 122608 115398
rect 153008 115954 153328 115986
rect 153008 115718 153050 115954
rect 153286 115718 153328 115954
rect 153008 115634 153328 115718
rect 153008 115398 153050 115634
rect 153286 115398 153328 115634
rect 153008 115366 153328 115398
rect 183728 115954 184048 115986
rect 183728 115718 183770 115954
rect 184006 115718 184048 115954
rect 183728 115634 184048 115718
rect 183728 115398 183770 115634
rect 184006 115398 184048 115634
rect 183728 115366 184048 115398
rect 214448 115954 214768 115986
rect 214448 115718 214490 115954
rect 214726 115718 214768 115954
rect 214448 115634 214768 115718
rect 214448 115398 214490 115634
rect 214726 115398 214768 115634
rect 214448 115366 214768 115398
rect 245168 115954 245488 115986
rect 245168 115718 245210 115954
rect 245446 115718 245488 115954
rect 245168 115634 245488 115718
rect 245168 115398 245210 115634
rect 245446 115398 245488 115634
rect 245168 115366 245488 115398
rect 275888 115954 276208 115986
rect 275888 115718 275930 115954
rect 276166 115718 276208 115954
rect 275888 115634 276208 115718
rect 275888 115398 275930 115634
rect 276166 115398 276208 115634
rect 275888 115366 276208 115398
rect 306608 115954 306928 115986
rect 306608 115718 306650 115954
rect 306886 115718 306928 115954
rect 306608 115634 306928 115718
rect 306608 115398 306650 115634
rect 306886 115398 306928 115634
rect 306608 115366 306928 115398
rect 337328 115954 337648 115986
rect 337328 115718 337370 115954
rect 337606 115718 337648 115954
rect 337328 115634 337648 115718
rect 337328 115398 337370 115634
rect 337606 115398 337648 115634
rect 337328 115366 337648 115398
rect 368048 115954 368368 115986
rect 368048 115718 368090 115954
rect 368326 115718 368368 115954
rect 368048 115634 368368 115718
rect 368048 115398 368090 115634
rect 368326 115398 368368 115634
rect 368048 115366 368368 115398
rect 398768 115954 399088 115986
rect 398768 115718 398810 115954
rect 399046 115718 399088 115954
rect 398768 115634 399088 115718
rect 398768 115398 398810 115634
rect 399046 115398 399088 115634
rect 398768 115366 399088 115398
rect 429488 115954 429808 115986
rect 429488 115718 429530 115954
rect 429766 115718 429808 115954
rect 429488 115634 429808 115718
rect 429488 115398 429530 115634
rect 429766 115398 429808 115634
rect 429488 115366 429808 115398
rect 460208 115954 460528 115986
rect 460208 115718 460250 115954
rect 460486 115718 460528 115954
rect 460208 115634 460528 115718
rect 460208 115398 460250 115634
rect 460486 115398 460528 115634
rect 460208 115366 460528 115398
rect 490928 115954 491248 115986
rect 490928 115718 490970 115954
rect 491206 115718 491248 115954
rect 490928 115634 491248 115718
rect 490928 115398 490970 115634
rect 491206 115398 491248 115634
rect 490928 115366 491248 115398
rect 76208 111454 76528 111486
rect 76208 111218 76250 111454
rect 76486 111218 76528 111454
rect 76208 111134 76528 111218
rect 76208 110898 76250 111134
rect 76486 110898 76528 111134
rect 76208 110866 76528 110898
rect 106928 111454 107248 111486
rect 106928 111218 106970 111454
rect 107206 111218 107248 111454
rect 106928 111134 107248 111218
rect 106928 110898 106970 111134
rect 107206 110898 107248 111134
rect 106928 110866 107248 110898
rect 137648 111454 137968 111486
rect 137648 111218 137690 111454
rect 137926 111218 137968 111454
rect 137648 111134 137968 111218
rect 137648 110898 137690 111134
rect 137926 110898 137968 111134
rect 137648 110866 137968 110898
rect 168368 111454 168688 111486
rect 168368 111218 168410 111454
rect 168646 111218 168688 111454
rect 168368 111134 168688 111218
rect 168368 110898 168410 111134
rect 168646 110898 168688 111134
rect 168368 110866 168688 110898
rect 199088 111454 199408 111486
rect 199088 111218 199130 111454
rect 199366 111218 199408 111454
rect 199088 111134 199408 111218
rect 199088 110898 199130 111134
rect 199366 110898 199408 111134
rect 199088 110866 199408 110898
rect 229808 111454 230128 111486
rect 229808 111218 229850 111454
rect 230086 111218 230128 111454
rect 229808 111134 230128 111218
rect 229808 110898 229850 111134
rect 230086 110898 230128 111134
rect 229808 110866 230128 110898
rect 260528 111454 260848 111486
rect 260528 111218 260570 111454
rect 260806 111218 260848 111454
rect 260528 111134 260848 111218
rect 260528 110898 260570 111134
rect 260806 110898 260848 111134
rect 260528 110866 260848 110898
rect 291248 111454 291568 111486
rect 291248 111218 291290 111454
rect 291526 111218 291568 111454
rect 291248 111134 291568 111218
rect 291248 110898 291290 111134
rect 291526 110898 291568 111134
rect 291248 110866 291568 110898
rect 321968 111454 322288 111486
rect 321968 111218 322010 111454
rect 322246 111218 322288 111454
rect 321968 111134 322288 111218
rect 321968 110898 322010 111134
rect 322246 110898 322288 111134
rect 321968 110866 322288 110898
rect 352688 111454 353008 111486
rect 352688 111218 352730 111454
rect 352966 111218 353008 111454
rect 352688 111134 353008 111218
rect 352688 110898 352730 111134
rect 352966 110898 353008 111134
rect 352688 110866 353008 110898
rect 383408 111454 383728 111486
rect 383408 111218 383450 111454
rect 383686 111218 383728 111454
rect 383408 111134 383728 111218
rect 383408 110898 383450 111134
rect 383686 110898 383728 111134
rect 383408 110866 383728 110898
rect 414128 111454 414448 111486
rect 414128 111218 414170 111454
rect 414406 111218 414448 111454
rect 414128 111134 414448 111218
rect 414128 110898 414170 111134
rect 414406 110898 414448 111134
rect 414128 110866 414448 110898
rect 444848 111454 445168 111486
rect 444848 111218 444890 111454
rect 445126 111218 445168 111454
rect 444848 111134 445168 111218
rect 444848 110898 444890 111134
rect 445126 110898 445168 111134
rect 444848 110866 445168 110898
rect 475568 111454 475888 111486
rect 475568 111218 475610 111454
rect 475846 111218 475888 111454
rect 475568 111134 475888 111218
rect 475568 110898 475610 111134
rect 475846 110898 475888 111134
rect 475568 110866 475888 110898
rect 506288 111454 506608 111486
rect 506288 111218 506330 111454
rect 506566 111218 506608 111454
rect 506288 111134 506608 111218
rect 506288 110898 506330 111134
rect 506566 110898 506608 111134
rect 506288 110866 506608 110898
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 91568 79954 91888 79986
rect 91568 79718 91610 79954
rect 91846 79718 91888 79954
rect 91568 79634 91888 79718
rect 91568 79398 91610 79634
rect 91846 79398 91888 79634
rect 91568 79366 91888 79398
rect 122288 79954 122608 79986
rect 122288 79718 122330 79954
rect 122566 79718 122608 79954
rect 122288 79634 122608 79718
rect 122288 79398 122330 79634
rect 122566 79398 122608 79634
rect 122288 79366 122608 79398
rect 153008 79954 153328 79986
rect 153008 79718 153050 79954
rect 153286 79718 153328 79954
rect 153008 79634 153328 79718
rect 153008 79398 153050 79634
rect 153286 79398 153328 79634
rect 153008 79366 153328 79398
rect 183728 79954 184048 79986
rect 183728 79718 183770 79954
rect 184006 79718 184048 79954
rect 183728 79634 184048 79718
rect 183728 79398 183770 79634
rect 184006 79398 184048 79634
rect 183728 79366 184048 79398
rect 214448 79954 214768 79986
rect 214448 79718 214490 79954
rect 214726 79718 214768 79954
rect 214448 79634 214768 79718
rect 214448 79398 214490 79634
rect 214726 79398 214768 79634
rect 214448 79366 214768 79398
rect 245168 79954 245488 79986
rect 245168 79718 245210 79954
rect 245446 79718 245488 79954
rect 245168 79634 245488 79718
rect 245168 79398 245210 79634
rect 245446 79398 245488 79634
rect 245168 79366 245488 79398
rect 275888 79954 276208 79986
rect 275888 79718 275930 79954
rect 276166 79718 276208 79954
rect 275888 79634 276208 79718
rect 275888 79398 275930 79634
rect 276166 79398 276208 79634
rect 275888 79366 276208 79398
rect 306608 79954 306928 79986
rect 306608 79718 306650 79954
rect 306886 79718 306928 79954
rect 306608 79634 306928 79718
rect 306608 79398 306650 79634
rect 306886 79398 306928 79634
rect 306608 79366 306928 79398
rect 337328 79954 337648 79986
rect 337328 79718 337370 79954
rect 337606 79718 337648 79954
rect 337328 79634 337648 79718
rect 337328 79398 337370 79634
rect 337606 79398 337648 79634
rect 337328 79366 337648 79398
rect 368048 79954 368368 79986
rect 368048 79718 368090 79954
rect 368326 79718 368368 79954
rect 368048 79634 368368 79718
rect 368048 79398 368090 79634
rect 368326 79398 368368 79634
rect 368048 79366 368368 79398
rect 398768 79954 399088 79986
rect 398768 79718 398810 79954
rect 399046 79718 399088 79954
rect 398768 79634 399088 79718
rect 398768 79398 398810 79634
rect 399046 79398 399088 79634
rect 398768 79366 399088 79398
rect 429488 79954 429808 79986
rect 429488 79718 429530 79954
rect 429766 79718 429808 79954
rect 429488 79634 429808 79718
rect 429488 79398 429530 79634
rect 429766 79398 429808 79634
rect 429488 79366 429808 79398
rect 460208 79954 460528 79986
rect 460208 79718 460250 79954
rect 460486 79718 460528 79954
rect 460208 79634 460528 79718
rect 460208 79398 460250 79634
rect 460486 79398 460528 79634
rect 460208 79366 460528 79398
rect 490928 79954 491248 79986
rect 490928 79718 490970 79954
rect 491206 79718 491248 79954
rect 490928 79634 491248 79718
rect 490928 79398 490970 79634
rect 491206 79398 491248 79634
rect 490928 79366 491248 79398
rect 76208 75454 76528 75486
rect 76208 75218 76250 75454
rect 76486 75218 76528 75454
rect 76208 75134 76528 75218
rect 76208 74898 76250 75134
rect 76486 74898 76528 75134
rect 76208 74866 76528 74898
rect 106928 75454 107248 75486
rect 106928 75218 106970 75454
rect 107206 75218 107248 75454
rect 106928 75134 107248 75218
rect 106928 74898 106970 75134
rect 107206 74898 107248 75134
rect 106928 74866 107248 74898
rect 137648 75454 137968 75486
rect 137648 75218 137690 75454
rect 137926 75218 137968 75454
rect 137648 75134 137968 75218
rect 137648 74898 137690 75134
rect 137926 74898 137968 75134
rect 137648 74866 137968 74898
rect 168368 75454 168688 75486
rect 168368 75218 168410 75454
rect 168646 75218 168688 75454
rect 168368 75134 168688 75218
rect 168368 74898 168410 75134
rect 168646 74898 168688 75134
rect 168368 74866 168688 74898
rect 199088 75454 199408 75486
rect 199088 75218 199130 75454
rect 199366 75218 199408 75454
rect 199088 75134 199408 75218
rect 199088 74898 199130 75134
rect 199366 74898 199408 75134
rect 199088 74866 199408 74898
rect 229808 75454 230128 75486
rect 229808 75218 229850 75454
rect 230086 75218 230128 75454
rect 229808 75134 230128 75218
rect 229808 74898 229850 75134
rect 230086 74898 230128 75134
rect 229808 74866 230128 74898
rect 260528 75454 260848 75486
rect 260528 75218 260570 75454
rect 260806 75218 260848 75454
rect 260528 75134 260848 75218
rect 260528 74898 260570 75134
rect 260806 74898 260848 75134
rect 260528 74866 260848 74898
rect 291248 75454 291568 75486
rect 291248 75218 291290 75454
rect 291526 75218 291568 75454
rect 291248 75134 291568 75218
rect 291248 74898 291290 75134
rect 291526 74898 291568 75134
rect 291248 74866 291568 74898
rect 321968 75454 322288 75486
rect 321968 75218 322010 75454
rect 322246 75218 322288 75454
rect 321968 75134 322288 75218
rect 321968 74898 322010 75134
rect 322246 74898 322288 75134
rect 321968 74866 322288 74898
rect 352688 75454 353008 75486
rect 352688 75218 352730 75454
rect 352966 75218 353008 75454
rect 352688 75134 353008 75218
rect 352688 74898 352730 75134
rect 352966 74898 353008 75134
rect 352688 74866 353008 74898
rect 383408 75454 383728 75486
rect 383408 75218 383450 75454
rect 383686 75218 383728 75454
rect 383408 75134 383728 75218
rect 383408 74898 383450 75134
rect 383686 74898 383728 75134
rect 383408 74866 383728 74898
rect 414128 75454 414448 75486
rect 414128 75218 414170 75454
rect 414406 75218 414448 75454
rect 414128 75134 414448 75218
rect 414128 74898 414170 75134
rect 414406 74898 414448 75134
rect 414128 74866 414448 74898
rect 444848 75454 445168 75486
rect 444848 75218 444890 75454
rect 445126 75218 445168 75454
rect 444848 75134 445168 75218
rect 444848 74898 444890 75134
rect 445126 74898 445168 75134
rect 444848 74866 445168 74898
rect 475568 75454 475888 75486
rect 475568 75218 475610 75454
rect 475846 75218 475888 75454
rect 475568 75134 475888 75218
rect 475568 74898 475610 75134
rect 475846 74898 475888 75134
rect 475568 74866 475888 74898
rect 506288 75454 506608 75486
rect 506288 75218 506330 75454
rect 506566 75218 506608 75454
rect 506288 75134 506608 75218
rect 506288 74898 506330 75134
rect 506566 74898 506608 75134
rect 506288 74866 506608 74898
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 39454 74414 70000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 43954 78914 70000
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 48454 83414 70000
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 52954 87914 70000
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 70000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 70000
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 70000
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 70000
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 70000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 70000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 70000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 70000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 70000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 70000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 70000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70000
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 39454 146414 70000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 70000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 70000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 70000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 70000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 70000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 70000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70000
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 70000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 70000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 70000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 70000
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 70000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 61954 204914 70000
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 66454 209414 70000
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 70000
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 39454 218414 70000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 43954 222914 70000
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 48454 227414 70000
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 52954 231914 70000
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 57454 236414 70000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 70000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 70000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 34954 249914 70000
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 39454 254414 70000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 43954 258914 70000
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 48454 263414 70000
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 52954 267914 70000
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 57454 272414 70000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 61954 276914 70000
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 66454 281414 70000
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 34954 285914 70000
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 39454 290414 70000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 43954 294914 70000
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 48454 299414 70000
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 52954 303914 70000
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 57454 308414 70000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 61954 312914 70000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 70000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 34954 321914 70000
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 39454 326414 70000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 43954 330914 70000
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 48454 335414 70000
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 52954 339914 70000
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 57454 344414 70000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 61954 348914 70000
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 66454 353414 70000
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 34954 357914 70000
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 39454 362414 70000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 43954 366914 70000
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 48454 371414 70000
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 52954 375914 70000
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 57454 380414 70000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 61954 384914 70000
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 66454 389414 70000
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 34954 393914 70000
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 39454 398414 70000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 43954 402914 70000
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 48454 407414 70000
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 52954 411914 70000
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 57454 416414 70000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 61954 420914 70000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 70000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 34954 429914 70000
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 39454 434414 70000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 43954 438914 70000
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 48454 443414 70000
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 52954 447914 70000
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 57454 452414 70000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 70000
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 66454 461414 70000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 34954 465914 70000
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 39454 470414 70000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 43954 474914 70000
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 48454 479414 70000
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 52954 483914 70000
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 57454 488414 70000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 61954 492914 70000
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 66454 497414 70000
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 34954 501914 70000
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 39454 506414 70000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 43954 510914 70000
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 580211 632364 580277 632365
rect 580211 632300 580212 632364
rect 580276 632300 580277 632364
rect 580211 632299 580277 632300
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 580214 139365 580274 632299
rect 580395 632092 580461 632093
rect 580395 632028 580396 632092
rect 580460 632028 580461 632092
rect 580395 632027 580461 632028
rect 580398 152693 580458 632027
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 580395 152692 580461 152693
rect 580395 152628 580396 152692
rect 580460 152628 580461 152692
rect 580395 152627 580461 152628
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 580211 139364 580277 139365
rect 580211 139300 580212 139364
rect 580276 139300 580277 139364
rect 580211 139299 580277 139300
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 91610 619718 91846 619954
rect 91610 619398 91846 619634
rect 122330 619718 122566 619954
rect 122330 619398 122566 619634
rect 153050 619718 153286 619954
rect 153050 619398 153286 619634
rect 183770 619718 184006 619954
rect 183770 619398 184006 619634
rect 214490 619718 214726 619954
rect 214490 619398 214726 619634
rect 245210 619718 245446 619954
rect 245210 619398 245446 619634
rect 275930 619718 276166 619954
rect 275930 619398 276166 619634
rect 306650 619718 306886 619954
rect 306650 619398 306886 619634
rect 337370 619718 337606 619954
rect 337370 619398 337606 619634
rect 368090 619718 368326 619954
rect 368090 619398 368326 619634
rect 398810 619718 399046 619954
rect 398810 619398 399046 619634
rect 429530 619718 429766 619954
rect 429530 619398 429766 619634
rect 460250 619718 460486 619954
rect 460250 619398 460486 619634
rect 490970 619718 491206 619954
rect 490970 619398 491206 619634
rect 76250 615218 76486 615454
rect 76250 614898 76486 615134
rect 106970 615218 107206 615454
rect 106970 614898 107206 615134
rect 137690 615218 137926 615454
rect 137690 614898 137926 615134
rect 168410 615218 168646 615454
rect 168410 614898 168646 615134
rect 199130 615218 199366 615454
rect 199130 614898 199366 615134
rect 229850 615218 230086 615454
rect 229850 614898 230086 615134
rect 260570 615218 260806 615454
rect 260570 614898 260806 615134
rect 291290 615218 291526 615454
rect 291290 614898 291526 615134
rect 322010 615218 322246 615454
rect 322010 614898 322246 615134
rect 352730 615218 352966 615454
rect 352730 614898 352966 615134
rect 383450 615218 383686 615454
rect 383450 614898 383686 615134
rect 414170 615218 414406 615454
rect 414170 614898 414406 615134
rect 444890 615218 445126 615454
rect 444890 614898 445126 615134
rect 475610 615218 475846 615454
rect 475610 614898 475846 615134
rect 506330 615218 506566 615454
rect 506330 614898 506566 615134
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 91610 583718 91846 583954
rect 91610 583398 91846 583634
rect 122330 583718 122566 583954
rect 122330 583398 122566 583634
rect 153050 583718 153286 583954
rect 153050 583398 153286 583634
rect 183770 583718 184006 583954
rect 183770 583398 184006 583634
rect 214490 583718 214726 583954
rect 214490 583398 214726 583634
rect 245210 583718 245446 583954
rect 245210 583398 245446 583634
rect 275930 583718 276166 583954
rect 275930 583398 276166 583634
rect 306650 583718 306886 583954
rect 306650 583398 306886 583634
rect 337370 583718 337606 583954
rect 337370 583398 337606 583634
rect 368090 583718 368326 583954
rect 368090 583398 368326 583634
rect 398810 583718 399046 583954
rect 398810 583398 399046 583634
rect 429530 583718 429766 583954
rect 429530 583398 429766 583634
rect 460250 583718 460486 583954
rect 460250 583398 460486 583634
rect 490970 583718 491206 583954
rect 490970 583398 491206 583634
rect 76250 579218 76486 579454
rect 76250 578898 76486 579134
rect 106970 579218 107206 579454
rect 106970 578898 107206 579134
rect 137690 579218 137926 579454
rect 137690 578898 137926 579134
rect 168410 579218 168646 579454
rect 168410 578898 168646 579134
rect 199130 579218 199366 579454
rect 199130 578898 199366 579134
rect 229850 579218 230086 579454
rect 229850 578898 230086 579134
rect 260570 579218 260806 579454
rect 260570 578898 260806 579134
rect 291290 579218 291526 579454
rect 291290 578898 291526 579134
rect 322010 579218 322246 579454
rect 322010 578898 322246 579134
rect 352730 579218 352966 579454
rect 352730 578898 352966 579134
rect 383450 579218 383686 579454
rect 383450 578898 383686 579134
rect 414170 579218 414406 579454
rect 414170 578898 414406 579134
rect 444890 579218 445126 579454
rect 444890 578898 445126 579134
rect 475610 579218 475846 579454
rect 475610 578898 475846 579134
rect 506330 579218 506566 579454
rect 506330 578898 506566 579134
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 91610 547718 91846 547954
rect 91610 547398 91846 547634
rect 122330 547718 122566 547954
rect 122330 547398 122566 547634
rect 153050 547718 153286 547954
rect 153050 547398 153286 547634
rect 183770 547718 184006 547954
rect 183770 547398 184006 547634
rect 214490 547718 214726 547954
rect 214490 547398 214726 547634
rect 245210 547718 245446 547954
rect 245210 547398 245446 547634
rect 275930 547718 276166 547954
rect 275930 547398 276166 547634
rect 306650 547718 306886 547954
rect 306650 547398 306886 547634
rect 337370 547718 337606 547954
rect 337370 547398 337606 547634
rect 368090 547718 368326 547954
rect 368090 547398 368326 547634
rect 398810 547718 399046 547954
rect 398810 547398 399046 547634
rect 429530 547718 429766 547954
rect 429530 547398 429766 547634
rect 460250 547718 460486 547954
rect 460250 547398 460486 547634
rect 490970 547718 491206 547954
rect 490970 547398 491206 547634
rect 76250 543218 76486 543454
rect 76250 542898 76486 543134
rect 106970 543218 107206 543454
rect 106970 542898 107206 543134
rect 137690 543218 137926 543454
rect 137690 542898 137926 543134
rect 168410 543218 168646 543454
rect 168410 542898 168646 543134
rect 199130 543218 199366 543454
rect 199130 542898 199366 543134
rect 229850 543218 230086 543454
rect 229850 542898 230086 543134
rect 260570 543218 260806 543454
rect 260570 542898 260806 543134
rect 291290 543218 291526 543454
rect 291290 542898 291526 543134
rect 322010 543218 322246 543454
rect 322010 542898 322246 543134
rect 352730 543218 352966 543454
rect 352730 542898 352966 543134
rect 383450 543218 383686 543454
rect 383450 542898 383686 543134
rect 414170 543218 414406 543454
rect 414170 542898 414406 543134
rect 444890 543218 445126 543454
rect 444890 542898 445126 543134
rect 475610 543218 475846 543454
rect 475610 542898 475846 543134
rect 506330 543218 506566 543454
rect 506330 542898 506566 543134
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 91610 511718 91846 511954
rect 91610 511398 91846 511634
rect 122330 511718 122566 511954
rect 122330 511398 122566 511634
rect 153050 511718 153286 511954
rect 153050 511398 153286 511634
rect 183770 511718 184006 511954
rect 183770 511398 184006 511634
rect 214490 511718 214726 511954
rect 214490 511398 214726 511634
rect 245210 511718 245446 511954
rect 245210 511398 245446 511634
rect 275930 511718 276166 511954
rect 275930 511398 276166 511634
rect 306650 511718 306886 511954
rect 306650 511398 306886 511634
rect 337370 511718 337606 511954
rect 337370 511398 337606 511634
rect 368090 511718 368326 511954
rect 368090 511398 368326 511634
rect 398810 511718 399046 511954
rect 398810 511398 399046 511634
rect 429530 511718 429766 511954
rect 429530 511398 429766 511634
rect 460250 511718 460486 511954
rect 460250 511398 460486 511634
rect 490970 511718 491206 511954
rect 490970 511398 491206 511634
rect 76250 507218 76486 507454
rect 76250 506898 76486 507134
rect 106970 507218 107206 507454
rect 106970 506898 107206 507134
rect 137690 507218 137926 507454
rect 137690 506898 137926 507134
rect 168410 507218 168646 507454
rect 168410 506898 168646 507134
rect 199130 507218 199366 507454
rect 199130 506898 199366 507134
rect 229850 507218 230086 507454
rect 229850 506898 230086 507134
rect 260570 507218 260806 507454
rect 260570 506898 260806 507134
rect 291290 507218 291526 507454
rect 291290 506898 291526 507134
rect 322010 507218 322246 507454
rect 322010 506898 322246 507134
rect 352730 507218 352966 507454
rect 352730 506898 352966 507134
rect 383450 507218 383686 507454
rect 383450 506898 383686 507134
rect 414170 507218 414406 507454
rect 414170 506898 414406 507134
rect 444890 507218 445126 507454
rect 444890 506898 445126 507134
rect 475610 507218 475846 507454
rect 475610 506898 475846 507134
rect 506330 507218 506566 507454
rect 506330 506898 506566 507134
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 91610 475718 91846 475954
rect 91610 475398 91846 475634
rect 122330 475718 122566 475954
rect 122330 475398 122566 475634
rect 153050 475718 153286 475954
rect 153050 475398 153286 475634
rect 183770 475718 184006 475954
rect 183770 475398 184006 475634
rect 214490 475718 214726 475954
rect 214490 475398 214726 475634
rect 245210 475718 245446 475954
rect 245210 475398 245446 475634
rect 275930 475718 276166 475954
rect 275930 475398 276166 475634
rect 306650 475718 306886 475954
rect 306650 475398 306886 475634
rect 337370 475718 337606 475954
rect 337370 475398 337606 475634
rect 368090 475718 368326 475954
rect 368090 475398 368326 475634
rect 398810 475718 399046 475954
rect 398810 475398 399046 475634
rect 429530 475718 429766 475954
rect 429530 475398 429766 475634
rect 460250 475718 460486 475954
rect 460250 475398 460486 475634
rect 490970 475718 491206 475954
rect 490970 475398 491206 475634
rect 76250 471218 76486 471454
rect 76250 470898 76486 471134
rect 106970 471218 107206 471454
rect 106970 470898 107206 471134
rect 137690 471218 137926 471454
rect 137690 470898 137926 471134
rect 168410 471218 168646 471454
rect 168410 470898 168646 471134
rect 199130 471218 199366 471454
rect 199130 470898 199366 471134
rect 229850 471218 230086 471454
rect 229850 470898 230086 471134
rect 260570 471218 260806 471454
rect 260570 470898 260806 471134
rect 291290 471218 291526 471454
rect 291290 470898 291526 471134
rect 322010 471218 322246 471454
rect 322010 470898 322246 471134
rect 352730 471218 352966 471454
rect 352730 470898 352966 471134
rect 383450 471218 383686 471454
rect 383450 470898 383686 471134
rect 414170 471218 414406 471454
rect 414170 470898 414406 471134
rect 444890 471218 445126 471454
rect 444890 470898 445126 471134
rect 475610 471218 475846 471454
rect 475610 470898 475846 471134
rect 506330 471218 506566 471454
rect 506330 470898 506566 471134
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 91610 439718 91846 439954
rect 91610 439398 91846 439634
rect 122330 439718 122566 439954
rect 122330 439398 122566 439634
rect 153050 439718 153286 439954
rect 153050 439398 153286 439634
rect 183770 439718 184006 439954
rect 183770 439398 184006 439634
rect 214490 439718 214726 439954
rect 214490 439398 214726 439634
rect 245210 439718 245446 439954
rect 245210 439398 245446 439634
rect 275930 439718 276166 439954
rect 275930 439398 276166 439634
rect 306650 439718 306886 439954
rect 306650 439398 306886 439634
rect 337370 439718 337606 439954
rect 337370 439398 337606 439634
rect 368090 439718 368326 439954
rect 368090 439398 368326 439634
rect 398810 439718 399046 439954
rect 398810 439398 399046 439634
rect 429530 439718 429766 439954
rect 429530 439398 429766 439634
rect 460250 439718 460486 439954
rect 460250 439398 460486 439634
rect 490970 439718 491206 439954
rect 490970 439398 491206 439634
rect 76250 435218 76486 435454
rect 76250 434898 76486 435134
rect 106970 435218 107206 435454
rect 106970 434898 107206 435134
rect 137690 435218 137926 435454
rect 137690 434898 137926 435134
rect 168410 435218 168646 435454
rect 168410 434898 168646 435134
rect 199130 435218 199366 435454
rect 199130 434898 199366 435134
rect 229850 435218 230086 435454
rect 229850 434898 230086 435134
rect 260570 435218 260806 435454
rect 260570 434898 260806 435134
rect 291290 435218 291526 435454
rect 291290 434898 291526 435134
rect 322010 435218 322246 435454
rect 322010 434898 322246 435134
rect 352730 435218 352966 435454
rect 352730 434898 352966 435134
rect 383450 435218 383686 435454
rect 383450 434898 383686 435134
rect 414170 435218 414406 435454
rect 414170 434898 414406 435134
rect 444890 435218 445126 435454
rect 444890 434898 445126 435134
rect 475610 435218 475846 435454
rect 475610 434898 475846 435134
rect 506330 435218 506566 435454
rect 506330 434898 506566 435134
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 91610 403718 91846 403954
rect 91610 403398 91846 403634
rect 122330 403718 122566 403954
rect 122330 403398 122566 403634
rect 153050 403718 153286 403954
rect 153050 403398 153286 403634
rect 183770 403718 184006 403954
rect 183770 403398 184006 403634
rect 214490 403718 214726 403954
rect 214490 403398 214726 403634
rect 245210 403718 245446 403954
rect 245210 403398 245446 403634
rect 275930 403718 276166 403954
rect 275930 403398 276166 403634
rect 306650 403718 306886 403954
rect 306650 403398 306886 403634
rect 337370 403718 337606 403954
rect 337370 403398 337606 403634
rect 368090 403718 368326 403954
rect 368090 403398 368326 403634
rect 398810 403718 399046 403954
rect 398810 403398 399046 403634
rect 429530 403718 429766 403954
rect 429530 403398 429766 403634
rect 460250 403718 460486 403954
rect 460250 403398 460486 403634
rect 490970 403718 491206 403954
rect 490970 403398 491206 403634
rect 76250 399218 76486 399454
rect 76250 398898 76486 399134
rect 106970 399218 107206 399454
rect 106970 398898 107206 399134
rect 137690 399218 137926 399454
rect 137690 398898 137926 399134
rect 168410 399218 168646 399454
rect 168410 398898 168646 399134
rect 199130 399218 199366 399454
rect 199130 398898 199366 399134
rect 229850 399218 230086 399454
rect 229850 398898 230086 399134
rect 260570 399218 260806 399454
rect 260570 398898 260806 399134
rect 291290 399218 291526 399454
rect 291290 398898 291526 399134
rect 322010 399218 322246 399454
rect 322010 398898 322246 399134
rect 352730 399218 352966 399454
rect 352730 398898 352966 399134
rect 383450 399218 383686 399454
rect 383450 398898 383686 399134
rect 414170 399218 414406 399454
rect 414170 398898 414406 399134
rect 444890 399218 445126 399454
rect 444890 398898 445126 399134
rect 475610 399218 475846 399454
rect 475610 398898 475846 399134
rect 506330 399218 506566 399454
rect 506330 398898 506566 399134
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 91610 367718 91846 367954
rect 91610 367398 91846 367634
rect 122330 367718 122566 367954
rect 122330 367398 122566 367634
rect 153050 367718 153286 367954
rect 153050 367398 153286 367634
rect 183770 367718 184006 367954
rect 183770 367398 184006 367634
rect 214490 367718 214726 367954
rect 214490 367398 214726 367634
rect 245210 367718 245446 367954
rect 245210 367398 245446 367634
rect 275930 367718 276166 367954
rect 275930 367398 276166 367634
rect 306650 367718 306886 367954
rect 306650 367398 306886 367634
rect 337370 367718 337606 367954
rect 337370 367398 337606 367634
rect 368090 367718 368326 367954
rect 368090 367398 368326 367634
rect 398810 367718 399046 367954
rect 398810 367398 399046 367634
rect 429530 367718 429766 367954
rect 429530 367398 429766 367634
rect 460250 367718 460486 367954
rect 460250 367398 460486 367634
rect 490970 367718 491206 367954
rect 490970 367398 491206 367634
rect 76250 363218 76486 363454
rect 76250 362898 76486 363134
rect 106970 363218 107206 363454
rect 106970 362898 107206 363134
rect 137690 363218 137926 363454
rect 137690 362898 137926 363134
rect 168410 363218 168646 363454
rect 168410 362898 168646 363134
rect 199130 363218 199366 363454
rect 199130 362898 199366 363134
rect 229850 363218 230086 363454
rect 229850 362898 230086 363134
rect 260570 363218 260806 363454
rect 260570 362898 260806 363134
rect 291290 363218 291526 363454
rect 291290 362898 291526 363134
rect 322010 363218 322246 363454
rect 322010 362898 322246 363134
rect 352730 363218 352966 363454
rect 352730 362898 352966 363134
rect 383450 363218 383686 363454
rect 383450 362898 383686 363134
rect 414170 363218 414406 363454
rect 414170 362898 414406 363134
rect 444890 363218 445126 363454
rect 444890 362898 445126 363134
rect 475610 363218 475846 363454
rect 475610 362898 475846 363134
rect 506330 363218 506566 363454
rect 506330 362898 506566 363134
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 91610 331718 91846 331954
rect 91610 331398 91846 331634
rect 122330 331718 122566 331954
rect 122330 331398 122566 331634
rect 153050 331718 153286 331954
rect 153050 331398 153286 331634
rect 183770 331718 184006 331954
rect 183770 331398 184006 331634
rect 214490 331718 214726 331954
rect 214490 331398 214726 331634
rect 245210 331718 245446 331954
rect 245210 331398 245446 331634
rect 275930 331718 276166 331954
rect 275930 331398 276166 331634
rect 306650 331718 306886 331954
rect 306650 331398 306886 331634
rect 337370 331718 337606 331954
rect 337370 331398 337606 331634
rect 368090 331718 368326 331954
rect 368090 331398 368326 331634
rect 398810 331718 399046 331954
rect 398810 331398 399046 331634
rect 429530 331718 429766 331954
rect 429530 331398 429766 331634
rect 460250 331718 460486 331954
rect 460250 331398 460486 331634
rect 490970 331718 491206 331954
rect 490970 331398 491206 331634
rect 76250 327218 76486 327454
rect 76250 326898 76486 327134
rect 106970 327218 107206 327454
rect 106970 326898 107206 327134
rect 137690 327218 137926 327454
rect 137690 326898 137926 327134
rect 168410 327218 168646 327454
rect 168410 326898 168646 327134
rect 199130 327218 199366 327454
rect 199130 326898 199366 327134
rect 229850 327218 230086 327454
rect 229850 326898 230086 327134
rect 260570 327218 260806 327454
rect 260570 326898 260806 327134
rect 291290 327218 291526 327454
rect 291290 326898 291526 327134
rect 322010 327218 322246 327454
rect 322010 326898 322246 327134
rect 352730 327218 352966 327454
rect 352730 326898 352966 327134
rect 383450 327218 383686 327454
rect 383450 326898 383686 327134
rect 414170 327218 414406 327454
rect 414170 326898 414406 327134
rect 444890 327218 445126 327454
rect 444890 326898 445126 327134
rect 475610 327218 475846 327454
rect 475610 326898 475846 327134
rect 506330 327218 506566 327454
rect 506330 326898 506566 327134
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 91610 295718 91846 295954
rect 91610 295398 91846 295634
rect 122330 295718 122566 295954
rect 122330 295398 122566 295634
rect 153050 295718 153286 295954
rect 153050 295398 153286 295634
rect 183770 295718 184006 295954
rect 183770 295398 184006 295634
rect 214490 295718 214726 295954
rect 214490 295398 214726 295634
rect 245210 295718 245446 295954
rect 245210 295398 245446 295634
rect 275930 295718 276166 295954
rect 275930 295398 276166 295634
rect 306650 295718 306886 295954
rect 306650 295398 306886 295634
rect 337370 295718 337606 295954
rect 337370 295398 337606 295634
rect 368090 295718 368326 295954
rect 368090 295398 368326 295634
rect 398810 295718 399046 295954
rect 398810 295398 399046 295634
rect 429530 295718 429766 295954
rect 429530 295398 429766 295634
rect 460250 295718 460486 295954
rect 460250 295398 460486 295634
rect 490970 295718 491206 295954
rect 490970 295398 491206 295634
rect 76250 291218 76486 291454
rect 76250 290898 76486 291134
rect 106970 291218 107206 291454
rect 106970 290898 107206 291134
rect 137690 291218 137926 291454
rect 137690 290898 137926 291134
rect 168410 291218 168646 291454
rect 168410 290898 168646 291134
rect 199130 291218 199366 291454
rect 199130 290898 199366 291134
rect 229850 291218 230086 291454
rect 229850 290898 230086 291134
rect 260570 291218 260806 291454
rect 260570 290898 260806 291134
rect 291290 291218 291526 291454
rect 291290 290898 291526 291134
rect 322010 291218 322246 291454
rect 322010 290898 322246 291134
rect 352730 291218 352966 291454
rect 352730 290898 352966 291134
rect 383450 291218 383686 291454
rect 383450 290898 383686 291134
rect 414170 291218 414406 291454
rect 414170 290898 414406 291134
rect 444890 291218 445126 291454
rect 444890 290898 445126 291134
rect 475610 291218 475846 291454
rect 475610 290898 475846 291134
rect 506330 291218 506566 291454
rect 506330 290898 506566 291134
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 91610 259718 91846 259954
rect 91610 259398 91846 259634
rect 122330 259718 122566 259954
rect 122330 259398 122566 259634
rect 153050 259718 153286 259954
rect 153050 259398 153286 259634
rect 183770 259718 184006 259954
rect 183770 259398 184006 259634
rect 214490 259718 214726 259954
rect 214490 259398 214726 259634
rect 245210 259718 245446 259954
rect 245210 259398 245446 259634
rect 275930 259718 276166 259954
rect 275930 259398 276166 259634
rect 306650 259718 306886 259954
rect 306650 259398 306886 259634
rect 337370 259718 337606 259954
rect 337370 259398 337606 259634
rect 368090 259718 368326 259954
rect 368090 259398 368326 259634
rect 398810 259718 399046 259954
rect 398810 259398 399046 259634
rect 429530 259718 429766 259954
rect 429530 259398 429766 259634
rect 460250 259718 460486 259954
rect 460250 259398 460486 259634
rect 490970 259718 491206 259954
rect 490970 259398 491206 259634
rect 76250 255218 76486 255454
rect 76250 254898 76486 255134
rect 106970 255218 107206 255454
rect 106970 254898 107206 255134
rect 137690 255218 137926 255454
rect 137690 254898 137926 255134
rect 168410 255218 168646 255454
rect 168410 254898 168646 255134
rect 199130 255218 199366 255454
rect 199130 254898 199366 255134
rect 229850 255218 230086 255454
rect 229850 254898 230086 255134
rect 260570 255218 260806 255454
rect 260570 254898 260806 255134
rect 291290 255218 291526 255454
rect 291290 254898 291526 255134
rect 322010 255218 322246 255454
rect 322010 254898 322246 255134
rect 352730 255218 352966 255454
rect 352730 254898 352966 255134
rect 383450 255218 383686 255454
rect 383450 254898 383686 255134
rect 414170 255218 414406 255454
rect 414170 254898 414406 255134
rect 444890 255218 445126 255454
rect 444890 254898 445126 255134
rect 475610 255218 475846 255454
rect 475610 254898 475846 255134
rect 506330 255218 506566 255454
rect 506330 254898 506566 255134
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 91610 223718 91846 223954
rect 91610 223398 91846 223634
rect 122330 223718 122566 223954
rect 122330 223398 122566 223634
rect 153050 223718 153286 223954
rect 153050 223398 153286 223634
rect 183770 223718 184006 223954
rect 183770 223398 184006 223634
rect 214490 223718 214726 223954
rect 214490 223398 214726 223634
rect 245210 223718 245446 223954
rect 245210 223398 245446 223634
rect 275930 223718 276166 223954
rect 275930 223398 276166 223634
rect 306650 223718 306886 223954
rect 306650 223398 306886 223634
rect 337370 223718 337606 223954
rect 337370 223398 337606 223634
rect 368090 223718 368326 223954
rect 368090 223398 368326 223634
rect 398810 223718 399046 223954
rect 398810 223398 399046 223634
rect 429530 223718 429766 223954
rect 429530 223398 429766 223634
rect 460250 223718 460486 223954
rect 460250 223398 460486 223634
rect 490970 223718 491206 223954
rect 490970 223398 491206 223634
rect 76250 219218 76486 219454
rect 76250 218898 76486 219134
rect 106970 219218 107206 219454
rect 106970 218898 107206 219134
rect 137690 219218 137926 219454
rect 137690 218898 137926 219134
rect 168410 219218 168646 219454
rect 168410 218898 168646 219134
rect 199130 219218 199366 219454
rect 199130 218898 199366 219134
rect 229850 219218 230086 219454
rect 229850 218898 230086 219134
rect 260570 219218 260806 219454
rect 260570 218898 260806 219134
rect 291290 219218 291526 219454
rect 291290 218898 291526 219134
rect 322010 219218 322246 219454
rect 322010 218898 322246 219134
rect 352730 219218 352966 219454
rect 352730 218898 352966 219134
rect 383450 219218 383686 219454
rect 383450 218898 383686 219134
rect 414170 219218 414406 219454
rect 414170 218898 414406 219134
rect 444890 219218 445126 219454
rect 444890 218898 445126 219134
rect 475610 219218 475846 219454
rect 475610 218898 475846 219134
rect 506330 219218 506566 219454
rect 506330 218898 506566 219134
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 91610 187718 91846 187954
rect 91610 187398 91846 187634
rect 122330 187718 122566 187954
rect 122330 187398 122566 187634
rect 153050 187718 153286 187954
rect 153050 187398 153286 187634
rect 183770 187718 184006 187954
rect 183770 187398 184006 187634
rect 214490 187718 214726 187954
rect 214490 187398 214726 187634
rect 245210 187718 245446 187954
rect 245210 187398 245446 187634
rect 275930 187718 276166 187954
rect 275930 187398 276166 187634
rect 306650 187718 306886 187954
rect 306650 187398 306886 187634
rect 337370 187718 337606 187954
rect 337370 187398 337606 187634
rect 368090 187718 368326 187954
rect 368090 187398 368326 187634
rect 398810 187718 399046 187954
rect 398810 187398 399046 187634
rect 429530 187718 429766 187954
rect 429530 187398 429766 187634
rect 460250 187718 460486 187954
rect 460250 187398 460486 187634
rect 490970 187718 491206 187954
rect 490970 187398 491206 187634
rect 76250 183218 76486 183454
rect 76250 182898 76486 183134
rect 106970 183218 107206 183454
rect 106970 182898 107206 183134
rect 137690 183218 137926 183454
rect 137690 182898 137926 183134
rect 168410 183218 168646 183454
rect 168410 182898 168646 183134
rect 199130 183218 199366 183454
rect 199130 182898 199366 183134
rect 229850 183218 230086 183454
rect 229850 182898 230086 183134
rect 260570 183218 260806 183454
rect 260570 182898 260806 183134
rect 291290 183218 291526 183454
rect 291290 182898 291526 183134
rect 322010 183218 322246 183454
rect 322010 182898 322246 183134
rect 352730 183218 352966 183454
rect 352730 182898 352966 183134
rect 383450 183218 383686 183454
rect 383450 182898 383686 183134
rect 414170 183218 414406 183454
rect 414170 182898 414406 183134
rect 444890 183218 445126 183454
rect 444890 182898 445126 183134
rect 475610 183218 475846 183454
rect 475610 182898 475846 183134
rect 506330 183218 506566 183454
rect 506330 182898 506566 183134
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 91610 151718 91846 151954
rect 91610 151398 91846 151634
rect 122330 151718 122566 151954
rect 122330 151398 122566 151634
rect 153050 151718 153286 151954
rect 153050 151398 153286 151634
rect 183770 151718 184006 151954
rect 183770 151398 184006 151634
rect 214490 151718 214726 151954
rect 214490 151398 214726 151634
rect 245210 151718 245446 151954
rect 245210 151398 245446 151634
rect 275930 151718 276166 151954
rect 275930 151398 276166 151634
rect 306650 151718 306886 151954
rect 306650 151398 306886 151634
rect 337370 151718 337606 151954
rect 337370 151398 337606 151634
rect 368090 151718 368326 151954
rect 368090 151398 368326 151634
rect 398810 151718 399046 151954
rect 398810 151398 399046 151634
rect 429530 151718 429766 151954
rect 429530 151398 429766 151634
rect 460250 151718 460486 151954
rect 460250 151398 460486 151634
rect 490970 151718 491206 151954
rect 490970 151398 491206 151634
rect 76250 147218 76486 147454
rect 76250 146898 76486 147134
rect 106970 147218 107206 147454
rect 106970 146898 107206 147134
rect 137690 147218 137926 147454
rect 137690 146898 137926 147134
rect 168410 147218 168646 147454
rect 168410 146898 168646 147134
rect 199130 147218 199366 147454
rect 199130 146898 199366 147134
rect 229850 147218 230086 147454
rect 229850 146898 230086 147134
rect 260570 147218 260806 147454
rect 260570 146898 260806 147134
rect 291290 147218 291526 147454
rect 291290 146898 291526 147134
rect 322010 147218 322246 147454
rect 322010 146898 322246 147134
rect 352730 147218 352966 147454
rect 352730 146898 352966 147134
rect 383450 147218 383686 147454
rect 383450 146898 383686 147134
rect 414170 147218 414406 147454
rect 414170 146898 414406 147134
rect 444890 147218 445126 147454
rect 444890 146898 445126 147134
rect 475610 147218 475846 147454
rect 475610 146898 475846 147134
rect 506330 147218 506566 147454
rect 506330 146898 506566 147134
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 91610 115718 91846 115954
rect 91610 115398 91846 115634
rect 122330 115718 122566 115954
rect 122330 115398 122566 115634
rect 153050 115718 153286 115954
rect 153050 115398 153286 115634
rect 183770 115718 184006 115954
rect 183770 115398 184006 115634
rect 214490 115718 214726 115954
rect 214490 115398 214726 115634
rect 245210 115718 245446 115954
rect 245210 115398 245446 115634
rect 275930 115718 276166 115954
rect 275930 115398 276166 115634
rect 306650 115718 306886 115954
rect 306650 115398 306886 115634
rect 337370 115718 337606 115954
rect 337370 115398 337606 115634
rect 368090 115718 368326 115954
rect 368090 115398 368326 115634
rect 398810 115718 399046 115954
rect 398810 115398 399046 115634
rect 429530 115718 429766 115954
rect 429530 115398 429766 115634
rect 460250 115718 460486 115954
rect 460250 115398 460486 115634
rect 490970 115718 491206 115954
rect 490970 115398 491206 115634
rect 76250 111218 76486 111454
rect 76250 110898 76486 111134
rect 106970 111218 107206 111454
rect 106970 110898 107206 111134
rect 137690 111218 137926 111454
rect 137690 110898 137926 111134
rect 168410 111218 168646 111454
rect 168410 110898 168646 111134
rect 199130 111218 199366 111454
rect 199130 110898 199366 111134
rect 229850 111218 230086 111454
rect 229850 110898 230086 111134
rect 260570 111218 260806 111454
rect 260570 110898 260806 111134
rect 291290 111218 291526 111454
rect 291290 110898 291526 111134
rect 322010 111218 322246 111454
rect 322010 110898 322246 111134
rect 352730 111218 352966 111454
rect 352730 110898 352966 111134
rect 383450 111218 383686 111454
rect 383450 110898 383686 111134
rect 414170 111218 414406 111454
rect 414170 110898 414406 111134
rect 444890 111218 445126 111454
rect 444890 110898 445126 111134
rect 475610 111218 475846 111454
rect 475610 110898 475846 111134
rect 506330 111218 506566 111454
rect 506330 110898 506566 111134
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 91610 79718 91846 79954
rect 91610 79398 91846 79634
rect 122330 79718 122566 79954
rect 122330 79398 122566 79634
rect 153050 79718 153286 79954
rect 153050 79398 153286 79634
rect 183770 79718 184006 79954
rect 183770 79398 184006 79634
rect 214490 79718 214726 79954
rect 214490 79398 214726 79634
rect 245210 79718 245446 79954
rect 245210 79398 245446 79634
rect 275930 79718 276166 79954
rect 275930 79398 276166 79634
rect 306650 79718 306886 79954
rect 306650 79398 306886 79634
rect 337370 79718 337606 79954
rect 337370 79398 337606 79634
rect 368090 79718 368326 79954
rect 368090 79398 368326 79634
rect 398810 79718 399046 79954
rect 398810 79398 399046 79634
rect 429530 79718 429766 79954
rect 429530 79398 429766 79634
rect 460250 79718 460486 79954
rect 460250 79398 460486 79634
rect 490970 79718 491206 79954
rect 490970 79398 491206 79634
rect 76250 75218 76486 75454
rect 76250 74898 76486 75134
rect 106970 75218 107206 75454
rect 106970 74898 107206 75134
rect 137690 75218 137926 75454
rect 137690 74898 137926 75134
rect 168410 75218 168646 75454
rect 168410 74898 168646 75134
rect 199130 75218 199366 75454
rect 199130 74898 199366 75134
rect 229850 75218 230086 75454
rect 229850 74898 230086 75134
rect 260570 75218 260806 75454
rect 260570 74898 260806 75134
rect 291290 75218 291526 75454
rect 291290 74898 291526 75134
rect 322010 75218 322246 75454
rect 322010 74898 322246 75134
rect 352730 75218 352966 75454
rect 352730 74898 352966 75134
rect 383450 75218 383686 75454
rect 383450 74898 383686 75134
rect 414170 75218 414406 75454
rect 414170 74898 414406 75134
rect 444890 75218 445126 75454
rect 444890 74898 445126 75134
rect 475610 75218 475846 75454
rect 475610 74898 475846 75134
rect 506330 75218 506566 75454
rect 506330 74898 506566 75134
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 91610 619954
rect 91846 619718 122330 619954
rect 122566 619718 153050 619954
rect 153286 619718 183770 619954
rect 184006 619718 214490 619954
rect 214726 619718 245210 619954
rect 245446 619718 275930 619954
rect 276166 619718 306650 619954
rect 306886 619718 337370 619954
rect 337606 619718 368090 619954
rect 368326 619718 398810 619954
rect 399046 619718 429530 619954
rect 429766 619718 460250 619954
rect 460486 619718 490970 619954
rect 491206 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 91610 619634
rect 91846 619398 122330 619634
rect 122566 619398 153050 619634
rect 153286 619398 183770 619634
rect 184006 619398 214490 619634
rect 214726 619398 245210 619634
rect 245446 619398 275930 619634
rect 276166 619398 306650 619634
rect 306886 619398 337370 619634
rect 337606 619398 368090 619634
rect 368326 619398 398810 619634
rect 399046 619398 429530 619634
rect 429766 619398 460250 619634
rect 460486 619398 490970 619634
rect 491206 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 76250 615454
rect 76486 615218 106970 615454
rect 107206 615218 137690 615454
rect 137926 615218 168410 615454
rect 168646 615218 199130 615454
rect 199366 615218 229850 615454
rect 230086 615218 260570 615454
rect 260806 615218 291290 615454
rect 291526 615218 322010 615454
rect 322246 615218 352730 615454
rect 352966 615218 383450 615454
rect 383686 615218 414170 615454
rect 414406 615218 444890 615454
rect 445126 615218 475610 615454
rect 475846 615218 506330 615454
rect 506566 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 76250 615134
rect 76486 614898 106970 615134
rect 107206 614898 137690 615134
rect 137926 614898 168410 615134
rect 168646 614898 199130 615134
rect 199366 614898 229850 615134
rect 230086 614898 260570 615134
rect 260806 614898 291290 615134
rect 291526 614898 322010 615134
rect 322246 614898 352730 615134
rect 352966 614898 383450 615134
rect 383686 614898 414170 615134
rect 414406 614898 444890 615134
rect 445126 614898 475610 615134
rect 475846 614898 506330 615134
rect 506566 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 91610 583954
rect 91846 583718 122330 583954
rect 122566 583718 153050 583954
rect 153286 583718 183770 583954
rect 184006 583718 214490 583954
rect 214726 583718 245210 583954
rect 245446 583718 275930 583954
rect 276166 583718 306650 583954
rect 306886 583718 337370 583954
rect 337606 583718 368090 583954
rect 368326 583718 398810 583954
rect 399046 583718 429530 583954
rect 429766 583718 460250 583954
rect 460486 583718 490970 583954
rect 491206 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 91610 583634
rect 91846 583398 122330 583634
rect 122566 583398 153050 583634
rect 153286 583398 183770 583634
rect 184006 583398 214490 583634
rect 214726 583398 245210 583634
rect 245446 583398 275930 583634
rect 276166 583398 306650 583634
rect 306886 583398 337370 583634
rect 337606 583398 368090 583634
rect 368326 583398 398810 583634
rect 399046 583398 429530 583634
rect 429766 583398 460250 583634
rect 460486 583398 490970 583634
rect 491206 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76250 579454
rect 76486 579218 106970 579454
rect 107206 579218 137690 579454
rect 137926 579218 168410 579454
rect 168646 579218 199130 579454
rect 199366 579218 229850 579454
rect 230086 579218 260570 579454
rect 260806 579218 291290 579454
rect 291526 579218 322010 579454
rect 322246 579218 352730 579454
rect 352966 579218 383450 579454
rect 383686 579218 414170 579454
rect 414406 579218 444890 579454
rect 445126 579218 475610 579454
rect 475846 579218 506330 579454
rect 506566 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76250 579134
rect 76486 578898 106970 579134
rect 107206 578898 137690 579134
rect 137926 578898 168410 579134
rect 168646 578898 199130 579134
rect 199366 578898 229850 579134
rect 230086 578898 260570 579134
rect 260806 578898 291290 579134
rect 291526 578898 322010 579134
rect 322246 578898 352730 579134
rect 352966 578898 383450 579134
rect 383686 578898 414170 579134
rect 414406 578898 444890 579134
rect 445126 578898 475610 579134
rect 475846 578898 506330 579134
rect 506566 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 91610 547954
rect 91846 547718 122330 547954
rect 122566 547718 153050 547954
rect 153286 547718 183770 547954
rect 184006 547718 214490 547954
rect 214726 547718 245210 547954
rect 245446 547718 275930 547954
rect 276166 547718 306650 547954
rect 306886 547718 337370 547954
rect 337606 547718 368090 547954
rect 368326 547718 398810 547954
rect 399046 547718 429530 547954
rect 429766 547718 460250 547954
rect 460486 547718 490970 547954
rect 491206 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 91610 547634
rect 91846 547398 122330 547634
rect 122566 547398 153050 547634
rect 153286 547398 183770 547634
rect 184006 547398 214490 547634
rect 214726 547398 245210 547634
rect 245446 547398 275930 547634
rect 276166 547398 306650 547634
rect 306886 547398 337370 547634
rect 337606 547398 368090 547634
rect 368326 547398 398810 547634
rect 399046 547398 429530 547634
rect 429766 547398 460250 547634
rect 460486 547398 490970 547634
rect 491206 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76250 543454
rect 76486 543218 106970 543454
rect 107206 543218 137690 543454
rect 137926 543218 168410 543454
rect 168646 543218 199130 543454
rect 199366 543218 229850 543454
rect 230086 543218 260570 543454
rect 260806 543218 291290 543454
rect 291526 543218 322010 543454
rect 322246 543218 352730 543454
rect 352966 543218 383450 543454
rect 383686 543218 414170 543454
rect 414406 543218 444890 543454
rect 445126 543218 475610 543454
rect 475846 543218 506330 543454
rect 506566 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76250 543134
rect 76486 542898 106970 543134
rect 107206 542898 137690 543134
rect 137926 542898 168410 543134
rect 168646 542898 199130 543134
rect 199366 542898 229850 543134
rect 230086 542898 260570 543134
rect 260806 542898 291290 543134
rect 291526 542898 322010 543134
rect 322246 542898 352730 543134
rect 352966 542898 383450 543134
rect 383686 542898 414170 543134
rect 414406 542898 444890 543134
rect 445126 542898 475610 543134
rect 475846 542898 506330 543134
rect 506566 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 91610 511954
rect 91846 511718 122330 511954
rect 122566 511718 153050 511954
rect 153286 511718 183770 511954
rect 184006 511718 214490 511954
rect 214726 511718 245210 511954
rect 245446 511718 275930 511954
rect 276166 511718 306650 511954
rect 306886 511718 337370 511954
rect 337606 511718 368090 511954
rect 368326 511718 398810 511954
rect 399046 511718 429530 511954
rect 429766 511718 460250 511954
rect 460486 511718 490970 511954
rect 491206 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 91610 511634
rect 91846 511398 122330 511634
rect 122566 511398 153050 511634
rect 153286 511398 183770 511634
rect 184006 511398 214490 511634
rect 214726 511398 245210 511634
rect 245446 511398 275930 511634
rect 276166 511398 306650 511634
rect 306886 511398 337370 511634
rect 337606 511398 368090 511634
rect 368326 511398 398810 511634
rect 399046 511398 429530 511634
rect 429766 511398 460250 511634
rect 460486 511398 490970 511634
rect 491206 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 76250 507454
rect 76486 507218 106970 507454
rect 107206 507218 137690 507454
rect 137926 507218 168410 507454
rect 168646 507218 199130 507454
rect 199366 507218 229850 507454
rect 230086 507218 260570 507454
rect 260806 507218 291290 507454
rect 291526 507218 322010 507454
rect 322246 507218 352730 507454
rect 352966 507218 383450 507454
rect 383686 507218 414170 507454
rect 414406 507218 444890 507454
rect 445126 507218 475610 507454
rect 475846 507218 506330 507454
rect 506566 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 76250 507134
rect 76486 506898 106970 507134
rect 107206 506898 137690 507134
rect 137926 506898 168410 507134
rect 168646 506898 199130 507134
rect 199366 506898 229850 507134
rect 230086 506898 260570 507134
rect 260806 506898 291290 507134
rect 291526 506898 322010 507134
rect 322246 506898 352730 507134
rect 352966 506898 383450 507134
rect 383686 506898 414170 507134
rect 414406 506898 444890 507134
rect 445126 506898 475610 507134
rect 475846 506898 506330 507134
rect 506566 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 91610 475954
rect 91846 475718 122330 475954
rect 122566 475718 153050 475954
rect 153286 475718 183770 475954
rect 184006 475718 214490 475954
rect 214726 475718 245210 475954
rect 245446 475718 275930 475954
rect 276166 475718 306650 475954
rect 306886 475718 337370 475954
rect 337606 475718 368090 475954
rect 368326 475718 398810 475954
rect 399046 475718 429530 475954
rect 429766 475718 460250 475954
rect 460486 475718 490970 475954
rect 491206 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 91610 475634
rect 91846 475398 122330 475634
rect 122566 475398 153050 475634
rect 153286 475398 183770 475634
rect 184006 475398 214490 475634
rect 214726 475398 245210 475634
rect 245446 475398 275930 475634
rect 276166 475398 306650 475634
rect 306886 475398 337370 475634
rect 337606 475398 368090 475634
rect 368326 475398 398810 475634
rect 399046 475398 429530 475634
rect 429766 475398 460250 475634
rect 460486 475398 490970 475634
rect 491206 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 76250 471454
rect 76486 471218 106970 471454
rect 107206 471218 137690 471454
rect 137926 471218 168410 471454
rect 168646 471218 199130 471454
rect 199366 471218 229850 471454
rect 230086 471218 260570 471454
rect 260806 471218 291290 471454
rect 291526 471218 322010 471454
rect 322246 471218 352730 471454
rect 352966 471218 383450 471454
rect 383686 471218 414170 471454
rect 414406 471218 444890 471454
rect 445126 471218 475610 471454
rect 475846 471218 506330 471454
rect 506566 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 76250 471134
rect 76486 470898 106970 471134
rect 107206 470898 137690 471134
rect 137926 470898 168410 471134
rect 168646 470898 199130 471134
rect 199366 470898 229850 471134
rect 230086 470898 260570 471134
rect 260806 470898 291290 471134
rect 291526 470898 322010 471134
rect 322246 470898 352730 471134
rect 352966 470898 383450 471134
rect 383686 470898 414170 471134
rect 414406 470898 444890 471134
rect 445126 470898 475610 471134
rect 475846 470898 506330 471134
rect 506566 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 91610 439954
rect 91846 439718 122330 439954
rect 122566 439718 153050 439954
rect 153286 439718 183770 439954
rect 184006 439718 214490 439954
rect 214726 439718 245210 439954
rect 245446 439718 275930 439954
rect 276166 439718 306650 439954
rect 306886 439718 337370 439954
rect 337606 439718 368090 439954
rect 368326 439718 398810 439954
rect 399046 439718 429530 439954
rect 429766 439718 460250 439954
rect 460486 439718 490970 439954
rect 491206 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 91610 439634
rect 91846 439398 122330 439634
rect 122566 439398 153050 439634
rect 153286 439398 183770 439634
rect 184006 439398 214490 439634
rect 214726 439398 245210 439634
rect 245446 439398 275930 439634
rect 276166 439398 306650 439634
rect 306886 439398 337370 439634
rect 337606 439398 368090 439634
rect 368326 439398 398810 439634
rect 399046 439398 429530 439634
rect 429766 439398 460250 439634
rect 460486 439398 490970 439634
rect 491206 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 76250 435454
rect 76486 435218 106970 435454
rect 107206 435218 137690 435454
rect 137926 435218 168410 435454
rect 168646 435218 199130 435454
rect 199366 435218 229850 435454
rect 230086 435218 260570 435454
rect 260806 435218 291290 435454
rect 291526 435218 322010 435454
rect 322246 435218 352730 435454
rect 352966 435218 383450 435454
rect 383686 435218 414170 435454
rect 414406 435218 444890 435454
rect 445126 435218 475610 435454
rect 475846 435218 506330 435454
rect 506566 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 76250 435134
rect 76486 434898 106970 435134
rect 107206 434898 137690 435134
rect 137926 434898 168410 435134
rect 168646 434898 199130 435134
rect 199366 434898 229850 435134
rect 230086 434898 260570 435134
rect 260806 434898 291290 435134
rect 291526 434898 322010 435134
rect 322246 434898 352730 435134
rect 352966 434898 383450 435134
rect 383686 434898 414170 435134
rect 414406 434898 444890 435134
rect 445126 434898 475610 435134
rect 475846 434898 506330 435134
rect 506566 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 91610 403954
rect 91846 403718 122330 403954
rect 122566 403718 153050 403954
rect 153286 403718 183770 403954
rect 184006 403718 214490 403954
rect 214726 403718 245210 403954
rect 245446 403718 275930 403954
rect 276166 403718 306650 403954
rect 306886 403718 337370 403954
rect 337606 403718 368090 403954
rect 368326 403718 398810 403954
rect 399046 403718 429530 403954
rect 429766 403718 460250 403954
rect 460486 403718 490970 403954
rect 491206 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 91610 403634
rect 91846 403398 122330 403634
rect 122566 403398 153050 403634
rect 153286 403398 183770 403634
rect 184006 403398 214490 403634
rect 214726 403398 245210 403634
rect 245446 403398 275930 403634
rect 276166 403398 306650 403634
rect 306886 403398 337370 403634
rect 337606 403398 368090 403634
rect 368326 403398 398810 403634
rect 399046 403398 429530 403634
rect 429766 403398 460250 403634
rect 460486 403398 490970 403634
rect 491206 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 76250 399454
rect 76486 399218 106970 399454
rect 107206 399218 137690 399454
rect 137926 399218 168410 399454
rect 168646 399218 199130 399454
rect 199366 399218 229850 399454
rect 230086 399218 260570 399454
rect 260806 399218 291290 399454
rect 291526 399218 322010 399454
rect 322246 399218 352730 399454
rect 352966 399218 383450 399454
rect 383686 399218 414170 399454
rect 414406 399218 444890 399454
rect 445126 399218 475610 399454
rect 475846 399218 506330 399454
rect 506566 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 76250 399134
rect 76486 398898 106970 399134
rect 107206 398898 137690 399134
rect 137926 398898 168410 399134
rect 168646 398898 199130 399134
rect 199366 398898 229850 399134
rect 230086 398898 260570 399134
rect 260806 398898 291290 399134
rect 291526 398898 322010 399134
rect 322246 398898 352730 399134
rect 352966 398898 383450 399134
rect 383686 398898 414170 399134
rect 414406 398898 444890 399134
rect 445126 398898 475610 399134
rect 475846 398898 506330 399134
rect 506566 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 91610 367954
rect 91846 367718 122330 367954
rect 122566 367718 153050 367954
rect 153286 367718 183770 367954
rect 184006 367718 214490 367954
rect 214726 367718 245210 367954
rect 245446 367718 275930 367954
rect 276166 367718 306650 367954
rect 306886 367718 337370 367954
rect 337606 367718 368090 367954
rect 368326 367718 398810 367954
rect 399046 367718 429530 367954
rect 429766 367718 460250 367954
rect 460486 367718 490970 367954
rect 491206 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 91610 367634
rect 91846 367398 122330 367634
rect 122566 367398 153050 367634
rect 153286 367398 183770 367634
rect 184006 367398 214490 367634
rect 214726 367398 245210 367634
rect 245446 367398 275930 367634
rect 276166 367398 306650 367634
rect 306886 367398 337370 367634
rect 337606 367398 368090 367634
rect 368326 367398 398810 367634
rect 399046 367398 429530 367634
rect 429766 367398 460250 367634
rect 460486 367398 490970 367634
rect 491206 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 76250 363454
rect 76486 363218 106970 363454
rect 107206 363218 137690 363454
rect 137926 363218 168410 363454
rect 168646 363218 199130 363454
rect 199366 363218 229850 363454
rect 230086 363218 260570 363454
rect 260806 363218 291290 363454
rect 291526 363218 322010 363454
rect 322246 363218 352730 363454
rect 352966 363218 383450 363454
rect 383686 363218 414170 363454
rect 414406 363218 444890 363454
rect 445126 363218 475610 363454
rect 475846 363218 506330 363454
rect 506566 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 76250 363134
rect 76486 362898 106970 363134
rect 107206 362898 137690 363134
rect 137926 362898 168410 363134
rect 168646 362898 199130 363134
rect 199366 362898 229850 363134
rect 230086 362898 260570 363134
rect 260806 362898 291290 363134
rect 291526 362898 322010 363134
rect 322246 362898 352730 363134
rect 352966 362898 383450 363134
rect 383686 362898 414170 363134
rect 414406 362898 444890 363134
rect 445126 362898 475610 363134
rect 475846 362898 506330 363134
rect 506566 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 91610 331954
rect 91846 331718 122330 331954
rect 122566 331718 153050 331954
rect 153286 331718 183770 331954
rect 184006 331718 214490 331954
rect 214726 331718 245210 331954
rect 245446 331718 275930 331954
rect 276166 331718 306650 331954
rect 306886 331718 337370 331954
rect 337606 331718 368090 331954
rect 368326 331718 398810 331954
rect 399046 331718 429530 331954
rect 429766 331718 460250 331954
rect 460486 331718 490970 331954
rect 491206 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 91610 331634
rect 91846 331398 122330 331634
rect 122566 331398 153050 331634
rect 153286 331398 183770 331634
rect 184006 331398 214490 331634
rect 214726 331398 245210 331634
rect 245446 331398 275930 331634
rect 276166 331398 306650 331634
rect 306886 331398 337370 331634
rect 337606 331398 368090 331634
rect 368326 331398 398810 331634
rect 399046 331398 429530 331634
rect 429766 331398 460250 331634
rect 460486 331398 490970 331634
rect 491206 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 76250 327454
rect 76486 327218 106970 327454
rect 107206 327218 137690 327454
rect 137926 327218 168410 327454
rect 168646 327218 199130 327454
rect 199366 327218 229850 327454
rect 230086 327218 260570 327454
rect 260806 327218 291290 327454
rect 291526 327218 322010 327454
rect 322246 327218 352730 327454
rect 352966 327218 383450 327454
rect 383686 327218 414170 327454
rect 414406 327218 444890 327454
rect 445126 327218 475610 327454
rect 475846 327218 506330 327454
rect 506566 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 76250 327134
rect 76486 326898 106970 327134
rect 107206 326898 137690 327134
rect 137926 326898 168410 327134
rect 168646 326898 199130 327134
rect 199366 326898 229850 327134
rect 230086 326898 260570 327134
rect 260806 326898 291290 327134
rect 291526 326898 322010 327134
rect 322246 326898 352730 327134
rect 352966 326898 383450 327134
rect 383686 326898 414170 327134
rect 414406 326898 444890 327134
rect 445126 326898 475610 327134
rect 475846 326898 506330 327134
rect 506566 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 91610 295954
rect 91846 295718 122330 295954
rect 122566 295718 153050 295954
rect 153286 295718 183770 295954
rect 184006 295718 214490 295954
rect 214726 295718 245210 295954
rect 245446 295718 275930 295954
rect 276166 295718 306650 295954
rect 306886 295718 337370 295954
rect 337606 295718 368090 295954
rect 368326 295718 398810 295954
rect 399046 295718 429530 295954
rect 429766 295718 460250 295954
rect 460486 295718 490970 295954
rect 491206 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 91610 295634
rect 91846 295398 122330 295634
rect 122566 295398 153050 295634
rect 153286 295398 183770 295634
rect 184006 295398 214490 295634
rect 214726 295398 245210 295634
rect 245446 295398 275930 295634
rect 276166 295398 306650 295634
rect 306886 295398 337370 295634
rect 337606 295398 368090 295634
rect 368326 295398 398810 295634
rect 399046 295398 429530 295634
rect 429766 295398 460250 295634
rect 460486 295398 490970 295634
rect 491206 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 76250 291454
rect 76486 291218 106970 291454
rect 107206 291218 137690 291454
rect 137926 291218 168410 291454
rect 168646 291218 199130 291454
rect 199366 291218 229850 291454
rect 230086 291218 260570 291454
rect 260806 291218 291290 291454
rect 291526 291218 322010 291454
rect 322246 291218 352730 291454
rect 352966 291218 383450 291454
rect 383686 291218 414170 291454
rect 414406 291218 444890 291454
rect 445126 291218 475610 291454
rect 475846 291218 506330 291454
rect 506566 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 76250 291134
rect 76486 290898 106970 291134
rect 107206 290898 137690 291134
rect 137926 290898 168410 291134
rect 168646 290898 199130 291134
rect 199366 290898 229850 291134
rect 230086 290898 260570 291134
rect 260806 290898 291290 291134
rect 291526 290898 322010 291134
rect 322246 290898 352730 291134
rect 352966 290898 383450 291134
rect 383686 290898 414170 291134
rect 414406 290898 444890 291134
rect 445126 290898 475610 291134
rect 475846 290898 506330 291134
rect 506566 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 91610 259954
rect 91846 259718 122330 259954
rect 122566 259718 153050 259954
rect 153286 259718 183770 259954
rect 184006 259718 214490 259954
rect 214726 259718 245210 259954
rect 245446 259718 275930 259954
rect 276166 259718 306650 259954
rect 306886 259718 337370 259954
rect 337606 259718 368090 259954
rect 368326 259718 398810 259954
rect 399046 259718 429530 259954
rect 429766 259718 460250 259954
rect 460486 259718 490970 259954
rect 491206 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 91610 259634
rect 91846 259398 122330 259634
rect 122566 259398 153050 259634
rect 153286 259398 183770 259634
rect 184006 259398 214490 259634
rect 214726 259398 245210 259634
rect 245446 259398 275930 259634
rect 276166 259398 306650 259634
rect 306886 259398 337370 259634
rect 337606 259398 368090 259634
rect 368326 259398 398810 259634
rect 399046 259398 429530 259634
rect 429766 259398 460250 259634
rect 460486 259398 490970 259634
rect 491206 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 76250 255454
rect 76486 255218 106970 255454
rect 107206 255218 137690 255454
rect 137926 255218 168410 255454
rect 168646 255218 199130 255454
rect 199366 255218 229850 255454
rect 230086 255218 260570 255454
rect 260806 255218 291290 255454
rect 291526 255218 322010 255454
rect 322246 255218 352730 255454
rect 352966 255218 383450 255454
rect 383686 255218 414170 255454
rect 414406 255218 444890 255454
rect 445126 255218 475610 255454
rect 475846 255218 506330 255454
rect 506566 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 76250 255134
rect 76486 254898 106970 255134
rect 107206 254898 137690 255134
rect 137926 254898 168410 255134
rect 168646 254898 199130 255134
rect 199366 254898 229850 255134
rect 230086 254898 260570 255134
rect 260806 254898 291290 255134
rect 291526 254898 322010 255134
rect 322246 254898 352730 255134
rect 352966 254898 383450 255134
rect 383686 254898 414170 255134
rect 414406 254898 444890 255134
rect 445126 254898 475610 255134
rect 475846 254898 506330 255134
rect 506566 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 91610 223954
rect 91846 223718 122330 223954
rect 122566 223718 153050 223954
rect 153286 223718 183770 223954
rect 184006 223718 214490 223954
rect 214726 223718 245210 223954
rect 245446 223718 275930 223954
rect 276166 223718 306650 223954
rect 306886 223718 337370 223954
rect 337606 223718 368090 223954
rect 368326 223718 398810 223954
rect 399046 223718 429530 223954
rect 429766 223718 460250 223954
rect 460486 223718 490970 223954
rect 491206 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 91610 223634
rect 91846 223398 122330 223634
rect 122566 223398 153050 223634
rect 153286 223398 183770 223634
rect 184006 223398 214490 223634
rect 214726 223398 245210 223634
rect 245446 223398 275930 223634
rect 276166 223398 306650 223634
rect 306886 223398 337370 223634
rect 337606 223398 368090 223634
rect 368326 223398 398810 223634
rect 399046 223398 429530 223634
rect 429766 223398 460250 223634
rect 460486 223398 490970 223634
rect 491206 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 76250 219454
rect 76486 219218 106970 219454
rect 107206 219218 137690 219454
rect 137926 219218 168410 219454
rect 168646 219218 199130 219454
rect 199366 219218 229850 219454
rect 230086 219218 260570 219454
rect 260806 219218 291290 219454
rect 291526 219218 322010 219454
rect 322246 219218 352730 219454
rect 352966 219218 383450 219454
rect 383686 219218 414170 219454
rect 414406 219218 444890 219454
rect 445126 219218 475610 219454
rect 475846 219218 506330 219454
rect 506566 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 76250 219134
rect 76486 218898 106970 219134
rect 107206 218898 137690 219134
rect 137926 218898 168410 219134
rect 168646 218898 199130 219134
rect 199366 218898 229850 219134
rect 230086 218898 260570 219134
rect 260806 218898 291290 219134
rect 291526 218898 322010 219134
rect 322246 218898 352730 219134
rect 352966 218898 383450 219134
rect 383686 218898 414170 219134
rect 414406 218898 444890 219134
rect 445126 218898 475610 219134
rect 475846 218898 506330 219134
rect 506566 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 91610 187954
rect 91846 187718 122330 187954
rect 122566 187718 153050 187954
rect 153286 187718 183770 187954
rect 184006 187718 214490 187954
rect 214726 187718 245210 187954
rect 245446 187718 275930 187954
rect 276166 187718 306650 187954
rect 306886 187718 337370 187954
rect 337606 187718 368090 187954
rect 368326 187718 398810 187954
rect 399046 187718 429530 187954
rect 429766 187718 460250 187954
rect 460486 187718 490970 187954
rect 491206 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 91610 187634
rect 91846 187398 122330 187634
rect 122566 187398 153050 187634
rect 153286 187398 183770 187634
rect 184006 187398 214490 187634
rect 214726 187398 245210 187634
rect 245446 187398 275930 187634
rect 276166 187398 306650 187634
rect 306886 187398 337370 187634
rect 337606 187398 368090 187634
rect 368326 187398 398810 187634
rect 399046 187398 429530 187634
rect 429766 187398 460250 187634
rect 460486 187398 490970 187634
rect 491206 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 76250 183454
rect 76486 183218 106970 183454
rect 107206 183218 137690 183454
rect 137926 183218 168410 183454
rect 168646 183218 199130 183454
rect 199366 183218 229850 183454
rect 230086 183218 260570 183454
rect 260806 183218 291290 183454
rect 291526 183218 322010 183454
rect 322246 183218 352730 183454
rect 352966 183218 383450 183454
rect 383686 183218 414170 183454
rect 414406 183218 444890 183454
rect 445126 183218 475610 183454
rect 475846 183218 506330 183454
rect 506566 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 76250 183134
rect 76486 182898 106970 183134
rect 107206 182898 137690 183134
rect 137926 182898 168410 183134
rect 168646 182898 199130 183134
rect 199366 182898 229850 183134
rect 230086 182898 260570 183134
rect 260806 182898 291290 183134
rect 291526 182898 322010 183134
rect 322246 182898 352730 183134
rect 352966 182898 383450 183134
rect 383686 182898 414170 183134
rect 414406 182898 444890 183134
rect 445126 182898 475610 183134
rect 475846 182898 506330 183134
rect 506566 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 91610 151954
rect 91846 151718 122330 151954
rect 122566 151718 153050 151954
rect 153286 151718 183770 151954
rect 184006 151718 214490 151954
rect 214726 151718 245210 151954
rect 245446 151718 275930 151954
rect 276166 151718 306650 151954
rect 306886 151718 337370 151954
rect 337606 151718 368090 151954
rect 368326 151718 398810 151954
rect 399046 151718 429530 151954
rect 429766 151718 460250 151954
rect 460486 151718 490970 151954
rect 491206 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 91610 151634
rect 91846 151398 122330 151634
rect 122566 151398 153050 151634
rect 153286 151398 183770 151634
rect 184006 151398 214490 151634
rect 214726 151398 245210 151634
rect 245446 151398 275930 151634
rect 276166 151398 306650 151634
rect 306886 151398 337370 151634
rect 337606 151398 368090 151634
rect 368326 151398 398810 151634
rect 399046 151398 429530 151634
rect 429766 151398 460250 151634
rect 460486 151398 490970 151634
rect 491206 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 76250 147454
rect 76486 147218 106970 147454
rect 107206 147218 137690 147454
rect 137926 147218 168410 147454
rect 168646 147218 199130 147454
rect 199366 147218 229850 147454
rect 230086 147218 260570 147454
rect 260806 147218 291290 147454
rect 291526 147218 322010 147454
rect 322246 147218 352730 147454
rect 352966 147218 383450 147454
rect 383686 147218 414170 147454
rect 414406 147218 444890 147454
rect 445126 147218 475610 147454
rect 475846 147218 506330 147454
rect 506566 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 76250 147134
rect 76486 146898 106970 147134
rect 107206 146898 137690 147134
rect 137926 146898 168410 147134
rect 168646 146898 199130 147134
rect 199366 146898 229850 147134
rect 230086 146898 260570 147134
rect 260806 146898 291290 147134
rect 291526 146898 322010 147134
rect 322246 146898 352730 147134
rect 352966 146898 383450 147134
rect 383686 146898 414170 147134
rect 414406 146898 444890 147134
rect 445126 146898 475610 147134
rect 475846 146898 506330 147134
rect 506566 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 91610 115954
rect 91846 115718 122330 115954
rect 122566 115718 153050 115954
rect 153286 115718 183770 115954
rect 184006 115718 214490 115954
rect 214726 115718 245210 115954
rect 245446 115718 275930 115954
rect 276166 115718 306650 115954
rect 306886 115718 337370 115954
rect 337606 115718 368090 115954
rect 368326 115718 398810 115954
rect 399046 115718 429530 115954
rect 429766 115718 460250 115954
rect 460486 115718 490970 115954
rect 491206 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 91610 115634
rect 91846 115398 122330 115634
rect 122566 115398 153050 115634
rect 153286 115398 183770 115634
rect 184006 115398 214490 115634
rect 214726 115398 245210 115634
rect 245446 115398 275930 115634
rect 276166 115398 306650 115634
rect 306886 115398 337370 115634
rect 337606 115398 368090 115634
rect 368326 115398 398810 115634
rect 399046 115398 429530 115634
rect 429766 115398 460250 115634
rect 460486 115398 490970 115634
rect 491206 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 76250 111454
rect 76486 111218 106970 111454
rect 107206 111218 137690 111454
rect 137926 111218 168410 111454
rect 168646 111218 199130 111454
rect 199366 111218 229850 111454
rect 230086 111218 260570 111454
rect 260806 111218 291290 111454
rect 291526 111218 322010 111454
rect 322246 111218 352730 111454
rect 352966 111218 383450 111454
rect 383686 111218 414170 111454
rect 414406 111218 444890 111454
rect 445126 111218 475610 111454
rect 475846 111218 506330 111454
rect 506566 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 76250 111134
rect 76486 110898 106970 111134
rect 107206 110898 137690 111134
rect 137926 110898 168410 111134
rect 168646 110898 199130 111134
rect 199366 110898 229850 111134
rect 230086 110898 260570 111134
rect 260806 110898 291290 111134
rect 291526 110898 322010 111134
rect 322246 110898 352730 111134
rect 352966 110898 383450 111134
rect 383686 110898 414170 111134
rect 414406 110898 444890 111134
rect 445126 110898 475610 111134
rect 475846 110898 506330 111134
rect 506566 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 91610 79954
rect 91846 79718 122330 79954
rect 122566 79718 153050 79954
rect 153286 79718 183770 79954
rect 184006 79718 214490 79954
rect 214726 79718 245210 79954
rect 245446 79718 275930 79954
rect 276166 79718 306650 79954
rect 306886 79718 337370 79954
rect 337606 79718 368090 79954
rect 368326 79718 398810 79954
rect 399046 79718 429530 79954
rect 429766 79718 460250 79954
rect 460486 79718 490970 79954
rect 491206 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 91610 79634
rect 91846 79398 122330 79634
rect 122566 79398 153050 79634
rect 153286 79398 183770 79634
rect 184006 79398 214490 79634
rect 214726 79398 245210 79634
rect 245446 79398 275930 79634
rect 276166 79398 306650 79634
rect 306886 79398 337370 79634
rect 337606 79398 368090 79634
rect 368326 79398 398810 79634
rect 399046 79398 429530 79634
rect 429766 79398 460250 79634
rect 460486 79398 490970 79634
rect 491206 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 76250 75454
rect 76486 75218 106970 75454
rect 107206 75218 137690 75454
rect 137926 75218 168410 75454
rect 168646 75218 199130 75454
rect 199366 75218 229850 75454
rect 230086 75218 260570 75454
rect 260806 75218 291290 75454
rect 291526 75218 322010 75454
rect 322246 75218 352730 75454
rect 352966 75218 383450 75454
rect 383686 75218 414170 75454
rect 414406 75218 444890 75454
rect 445126 75218 475610 75454
rect 475846 75218 506330 75454
rect 506566 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 76250 75134
rect 76486 74898 106970 75134
rect 107206 74898 137690 75134
rect 137926 74898 168410 75134
rect 168646 74898 199130 75134
rect 199366 74898 229850 75134
rect 230086 74898 260570 75134
rect 260806 74898 291290 75134
rect 291526 74898 322010 75134
rect 322246 74898 352730 75134
rect 352966 74898 383450 75134
rect 383686 74898 414170 75134
rect 414406 74898 444890 75134
rect 445126 74898 475610 75134
rect 475846 74898 506330 75134
rect 506566 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use trainable_nn  mprj
timestamp 0
transform 1 0 72000 0 1 72000
box 1066 0 439011 560000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 634000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 634000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 634000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 634000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 634000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 634000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 634000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 634000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 634000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 634000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 634000 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 634000 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 70000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 634000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 634000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 634000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 634000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 634000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 634000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 634000 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 634000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 634000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 634000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 634000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 634000 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 70000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 634000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 634000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 634000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 634000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 634000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 634000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 634000 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 634000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 634000 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 634000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 634000 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 634000 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 70000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 634000 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 634000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 634000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 634000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 634000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 634000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 634000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 634000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 634000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 634000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 634000 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 634000 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 70000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 634000 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 634000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 634000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 634000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 634000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 634000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 634000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 634000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 634000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 634000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 634000 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 634000 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 70000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 634000 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 634000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 634000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 634000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 634000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 634000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 634000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 634000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 634000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 634000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 634000 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 634000 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 70000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 634000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 634000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 634000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 634000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 634000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 634000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 634000 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 634000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 634000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 634000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 634000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 634000 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 634000 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 70000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 634000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 634000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 634000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 634000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 634000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 634000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 634000 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 634000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 634000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 634000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 634000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 634000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 70000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 634000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
