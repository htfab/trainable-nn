magic
tech sky130B
magscale 1 2
timestamp 1663048280
<< nwell >>
rect 1066 557317 438878 557638
rect 1066 556229 438878 556795
rect 1066 555141 438878 555707
rect 1066 554053 438878 554619
rect 1066 552965 438878 553531
rect 1066 551877 438878 552443
rect 1066 550789 438878 551355
rect 1066 549701 438878 550267
rect 1066 548613 438878 549179
rect 1066 547525 438878 548091
rect 1066 546437 438878 547003
rect 1066 545349 438878 545915
rect 1066 544261 438878 544827
rect 1066 543173 438878 543739
rect 1066 542085 438878 542651
rect 1066 540997 438878 541563
rect 1066 539909 438878 540475
rect 1066 538821 438878 539387
rect 1066 537733 438878 538299
rect 1066 536645 438878 537211
rect 1066 535557 438878 536123
rect 1066 534469 438878 535035
rect 1066 533381 438878 533947
rect 1066 532293 438878 532859
rect 1066 531205 438878 531771
rect 1066 530117 438878 530683
rect 1066 529029 438878 529595
rect 1066 527941 438878 528507
rect 1066 526853 438878 527419
rect 1066 525765 438878 526331
rect 1066 524677 438878 525243
rect 1066 523589 438878 524155
rect 1066 522501 438878 523067
rect 1066 521413 438878 521979
rect 1066 520325 438878 520891
rect 1066 519237 438878 519803
rect 1066 518149 438878 518715
rect 1066 517061 438878 517627
rect 1066 515973 438878 516539
rect 1066 514885 438878 515451
rect 1066 513797 438878 514363
rect 1066 512709 438878 513275
rect 1066 511621 438878 512187
rect 1066 510533 438878 511099
rect 1066 509445 438878 510011
rect 1066 508357 438878 508923
rect 1066 507269 438878 507835
rect 1066 506181 438878 506747
rect 1066 505093 438878 505659
rect 1066 504005 438878 504571
rect 1066 502917 438878 503483
rect 1066 501829 438878 502395
rect 1066 500741 438878 501307
rect 1066 499653 438878 500219
rect 1066 498565 438878 499131
rect 1066 497477 438878 498043
rect 1066 496389 438878 496955
rect 1066 495301 438878 495867
rect 1066 494213 438878 494779
rect 1066 493125 438878 493691
rect 1066 492037 438878 492603
rect 1066 490949 438878 491515
rect 1066 489861 438878 490427
rect 1066 488773 438878 489339
rect 1066 487685 438878 488251
rect 1066 486597 438878 487163
rect 1066 485509 438878 486075
rect 1066 484421 438878 484987
rect 1066 483333 438878 483899
rect 1066 482245 438878 482811
rect 1066 481157 438878 481723
rect 1066 480069 438878 480635
rect 1066 478981 438878 479547
rect 1066 477893 438878 478459
rect 1066 476805 438878 477371
rect 1066 475717 438878 476283
rect 1066 474629 438878 475195
rect 1066 473541 438878 474107
rect 1066 472453 438878 473019
rect 1066 471365 438878 471931
rect 1066 470277 438878 470843
rect 1066 469189 438878 469755
rect 1066 468101 438878 468667
rect 1066 467013 438878 467579
rect 1066 465925 438878 466491
rect 1066 464837 438878 465403
rect 1066 463749 438878 464315
rect 1066 462661 438878 463227
rect 1066 461573 438878 462139
rect 1066 460485 438878 461051
rect 1066 459397 438878 459963
rect 1066 458309 438878 458875
rect 1066 457221 438878 457787
rect 1066 456133 438878 456699
rect 1066 455045 438878 455611
rect 1066 453957 438878 454523
rect 1066 452869 438878 453435
rect 1066 451781 438878 452347
rect 1066 450693 438878 451259
rect 1066 449605 438878 450171
rect 1066 448517 438878 449083
rect 1066 447429 438878 447995
rect 1066 446341 438878 446907
rect 1066 445253 438878 445819
rect 1066 444165 438878 444731
rect 1066 443077 438878 443643
rect 1066 441989 438878 442555
rect 1066 440901 438878 441467
rect 1066 439813 438878 440379
rect 1066 438725 438878 439291
rect 1066 437637 438878 438203
rect 1066 436549 438878 437115
rect 1066 435461 438878 436027
rect 1066 434373 438878 434939
rect 1066 433285 438878 433851
rect 1066 432197 438878 432763
rect 1066 431109 438878 431675
rect 1066 430021 438878 430587
rect 1066 428933 438878 429499
rect 1066 427845 438878 428411
rect 1066 426757 438878 427323
rect 1066 425669 438878 426235
rect 1066 424581 438878 425147
rect 1066 423493 438878 424059
rect 1066 422405 438878 422971
rect 1066 421317 438878 421883
rect 1066 420229 438878 420795
rect 1066 419141 438878 419707
rect 1066 418053 438878 418619
rect 1066 416965 438878 417531
rect 1066 415877 438878 416443
rect 1066 414789 438878 415355
rect 1066 413701 438878 414267
rect 1066 412613 438878 413179
rect 1066 411525 438878 412091
rect 1066 410437 438878 411003
rect 1066 409349 438878 409915
rect 1066 408261 438878 408827
rect 1066 407173 438878 407739
rect 1066 406085 438878 406651
rect 1066 404997 438878 405563
rect 1066 403909 438878 404475
rect 1066 402821 438878 403387
rect 1066 401733 438878 402299
rect 1066 400645 438878 401211
rect 1066 399557 438878 400123
rect 1066 398469 438878 399035
rect 1066 397381 438878 397947
rect 1066 396293 438878 396859
rect 1066 395205 438878 395771
rect 1066 394117 438878 394683
rect 1066 393029 438878 393595
rect 1066 391941 438878 392507
rect 1066 390853 438878 391419
rect 1066 389765 438878 390331
rect 1066 388677 438878 389243
rect 1066 387589 438878 388155
rect 1066 386501 438878 387067
rect 1066 385413 438878 385979
rect 1066 384325 438878 384891
rect 1066 383237 438878 383803
rect 1066 382149 438878 382715
rect 1066 381061 438878 381627
rect 1066 379973 438878 380539
rect 1066 378885 438878 379451
rect 1066 377797 438878 378363
rect 1066 376709 438878 377275
rect 1066 375621 438878 376187
rect 1066 374533 438878 375099
rect 1066 373445 438878 374011
rect 1066 372357 438878 372923
rect 1066 371269 438878 371835
rect 1066 370181 438878 370747
rect 1066 369093 438878 369659
rect 1066 368005 438878 368571
rect 1066 366917 438878 367483
rect 1066 365829 438878 366395
rect 1066 364741 438878 365307
rect 1066 363653 438878 364219
rect 1066 362565 438878 363131
rect 1066 361477 438878 362043
rect 1066 360389 438878 360955
rect 1066 359301 438878 359867
rect 1066 358213 438878 358779
rect 1066 357125 438878 357691
rect 1066 356037 438878 356603
rect 1066 354949 438878 355515
rect 1066 353861 438878 354427
rect 1066 352773 438878 353339
rect 1066 351685 438878 352251
rect 1066 350597 438878 351163
rect 1066 349509 438878 350075
rect 1066 348421 438878 348987
rect 1066 347333 438878 347899
rect 1066 346245 438878 346811
rect 1066 345157 438878 345723
rect 1066 344069 438878 344635
rect 1066 342981 438878 343547
rect 1066 341893 438878 342459
rect 1066 340805 438878 341371
rect 1066 339717 438878 340283
rect 1066 338629 438878 339195
rect 1066 337541 438878 338107
rect 1066 336453 438878 337019
rect 1066 335365 438878 335931
rect 1066 334277 438878 334843
rect 1066 333189 438878 333755
rect 1066 332101 438878 332667
rect 1066 331013 438878 331579
rect 1066 329925 438878 330491
rect 1066 328837 438878 329403
rect 1066 327749 438878 328315
rect 1066 326661 438878 327227
rect 1066 325573 438878 326139
rect 1066 324485 438878 325051
rect 1066 323397 438878 323963
rect 1066 322309 438878 322875
rect 1066 321221 438878 321787
rect 1066 320133 438878 320699
rect 1066 319045 438878 319611
rect 1066 317957 438878 318523
rect 1066 316869 438878 317435
rect 1066 315781 438878 316347
rect 1066 314693 438878 315259
rect 1066 313605 438878 314171
rect 1066 312517 438878 313083
rect 1066 311429 438878 311995
rect 1066 310341 438878 310907
rect 1066 309253 438878 309819
rect 1066 308165 438878 308731
rect 1066 307077 438878 307643
rect 1066 305989 438878 306555
rect 1066 304901 438878 305467
rect 1066 303813 438878 304379
rect 1066 302725 438878 303291
rect 1066 301637 438878 302203
rect 1066 300549 438878 301115
rect 1066 299461 438878 300027
rect 1066 298373 438878 298939
rect 1066 297285 438878 297851
rect 1066 296197 438878 296763
rect 1066 295109 438878 295675
rect 1066 294021 438878 294587
rect 1066 292933 438878 293499
rect 1066 291845 438878 292411
rect 1066 290757 438878 291323
rect 1066 289669 438878 290235
rect 1066 288581 438878 289147
rect 1066 287493 438878 288059
rect 1066 286405 438878 286971
rect 1066 285317 438878 285883
rect 1066 284229 438878 284795
rect 1066 283141 438878 283707
rect 1066 282053 438878 282619
rect 1066 280965 438878 281531
rect 1066 279877 438878 280443
rect 1066 278789 438878 279355
rect 1066 277701 438878 278267
rect 1066 276613 438878 277179
rect 1066 275525 438878 276091
rect 1066 274437 438878 275003
rect 1066 273349 438878 273915
rect 1066 272261 438878 272827
rect 1066 271173 438878 271739
rect 1066 270085 438878 270651
rect 1066 268997 438878 269563
rect 1066 267909 438878 268475
rect 1066 266821 438878 267387
rect 1066 265733 438878 266299
rect 1066 264645 438878 265211
rect 1066 263557 438878 264123
rect 1066 262469 438878 263035
rect 1066 261381 438878 261947
rect 1066 260293 438878 260859
rect 1066 259205 438878 259771
rect 1066 258117 438878 258683
rect 1066 257029 438878 257595
rect 1066 255941 438878 256507
rect 1066 254853 438878 255419
rect 1066 253765 438878 254331
rect 1066 252677 438878 253243
rect 1066 251589 438878 252155
rect 1066 250501 438878 251067
rect 1066 249413 438878 249979
rect 1066 248325 438878 248891
rect 1066 247237 438878 247803
rect 1066 246149 438878 246715
rect 1066 245061 438878 245627
rect 1066 243973 438878 244539
rect 1066 242885 438878 243451
rect 1066 241797 438878 242363
rect 1066 240709 438878 241275
rect 1066 239621 438878 240187
rect 1066 238533 438878 239099
rect 1066 237445 438878 238011
rect 1066 236357 438878 236923
rect 1066 235269 438878 235835
rect 1066 234181 438878 234747
rect 1066 233093 438878 233659
rect 1066 232005 438878 232571
rect 1066 230917 438878 231483
rect 1066 229829 438878 230395
rect 1066 228741 438878 229307
rect 1066 227653 438878 228219
rect 1066 226565 438878 227131
rect 1066 225477 438878 226043
rect 1066 224389 438878 224955
rect 1066 223301 438878 223867
rect 1066 222213 438878 222779
rect 1066 221125 438878 221691
rect 1066 220037 438878 220603
rect 1066 218949 438878 219515
rect 1066 217861 438878 218427
rect 1066 216773 438878 217339
rect 1066 215685 438878 216251
rect 1066 214597 438878 215163
rect 1066 213509 438878 214075
rect 1066 212421 438878 212987
rect 1066 211333 438878 211899
rect 1066 210245 438878 210811
rect 1066 209157 438878 209723
rect 1066 208069 438878 208635
rect 1066 206981 438878 207547
rect 1066 205893 438878 206459
rect 1066 204805 438878 205371
rect 1066 203717 438878 204283
rect 1066 202629 438878 203195
rect 1066 201541 438878 202107
rect 1066 200453 438878 201019
rect 1066 199365 438878 199931
rect 1066 198277 438878 198843
rect 1066 197189 438878 197755
rect 1066 196101 438878 196667
rect 1066 195013 438878 195579
rect 1066 193925 438878 194491
rect 1066 192837 438878 193403
rect 1066 191749 438878 192315
rect 1066 190661 438878 191227
rect 1066 189573 438878 190139
rect 1066 188485 438878 189051
rect 1066 187397 438878 187963
rect 1066 186309 438878 186875
rect 1066 185221 438878 185787
rect 1066 184133 438878 184699
rect 1066 183045 438878 183611
rect 1066 181957 438878 182523
rect 1066 180869 438878 181435
rect 1066 179781 438878 180347
rect 1066 178693 438878 179259
rect 1066 177605 438878 178171
rect 1066 176517 438878 177083
rect 1066 175429 438878 175995
rect 1066 174341 438878 174907
rect 1066 173253 438878 173819
rect 1066 172165 438878 172731
rect 1066 171077 438878 171643
rect 1066 169989 438878 170555
rect 1066 168901 438878 169467
rect 1066 167813 438878 168379
rect 1066 166725 438878 167291
rect 1066 165637 438878 166203
rect 1066 164549 438878 165115
rect 1066 163461 438878 164027
rect 1066 162373 438878 162939
rect 1066 161285 438878 161851
rect 1066 160197 438878 160763
rect 1066 159109 438878 159675
rect 1066 158021 438878 158587
rect 1066 156933 438878 157499
rect 1066 155845 438878 156411
rect 1066 154757 438878 155323
rect 1066 153669 438878 154235
rect 1066 152581 438878 153147
rect 1066 151493 438878 152059
rect 1066 150405 438878 150971
rect 1066 149317 438878 149883
rect 1066 148229 438878 148795
rect 1066 147141 438878 147707
rect 1066 146053 438878 146619
rect 1066 144965 438878 145531
rect 1066 143877 438878 144443
rect 1066 142789 438878 143355
rect 1066 141701 438878 142267
rect 1066 140613 438878 141179
rect 1066 139525 438878 140091
rect 1066 138437 438878 139003
rect 1066 137349 438878 137915
rect 1066 136261 438878 136827
rect 1066 135173 438878 135739
rect 1066 134085 438878 134651
rect 1066 132997 438878 133563
rect 1066 131909 438878 132475
rect 1066 130821 438878 131387
rect 1066 129733 438878 130299
rect 1066 128645 438878 129211
rect 1066 127557 438878 128123
rect 1066 126469 438878 127035
rect 1066 125381 438878 125947
rect 1066 124293 438878 124859
rect 1066 123205 438878 123771
rect 1066 122117 438878 122683
rect 1066 121029 438878 121595
rect 1066 119941 438878 120507
rect 1066 118853 438878 119419
rect 1066 117765 438878 118331
rect 1066 116677 438878 117243
rect 1066 115589 438878 116155
rect 1066 114501 438878 115067
rect 1066 113413 438878 113979
rect 1066 112325 438878 112891
rect 1066 111237 438878 111803
rect 1066 110149 438878 110715
rect 1066 109061 438878 109627
rect 1066 107973 438878 108539
rect 1066 106885 438878 107451
rect 1066 105797 438878 106363
rect 1066 104709 438878 105275
rect 1066 103621 438878 104187
rect 1066 102533 438878 103099
rect 1066 101445 438878 102011
rect 1066 100357 438878 100923
rect 1066 99269 438878 99835
rect 1066 98181 438878 98747
rect 1066 97093 438878 97659
rect 1066 96005 438878 96571
rect 1066 94917 438878 95483
rect 1066 93829 438878 94395
rect 1066 92741 438878 93307
rect 1066 91653 438878 92219
rect 1066 90565 438878 91131
rect 1066 89477 438878 90043
rect 1066 88389 438878 88955
rect 1066 87301 438878 87867
rect 1066 86213 438878 86779
rect 1066 85125 438878 85691
rect 1066 84037 438878 84603
rect 1066 82949 438878 83515
rect 1066 81861 438878 82427
rect 1066 80773 438878 81339
rect 1066 79685 438878 80251
rect 1066 78597 438878 79163
rect 1066 77509 438878 78075
rect 1066 76421 438878 76987
rect 1066 75333 438878 75899
rect 1066 74245 438878 74811
rect 1066 73157 438878 73723
rect 1066 72069 438878 72635
rect 1066 70981 438878 71547
rect 1066 69893 438878 70459
rect 1066 68805 438878 69371
rect 1066 67717 438878 68283
rect 1066 66629 438878 67195
rect 1066 65541 438878 66107
rect 1066 64453 438878 65019
rect 1066 63365 438878 63931
rect 1066 62277 438878 62843
rect 1066 61189 438878 61755
rect 1066 60101 438878 60667
rect 1066 59013 438878 59579
rect 1066 57925 438878 58491
rect 1066 56837 438878 57403
rect 1066 55749 438878 56315
rect 1066 54661 438878 55227
rect 1066 53573 438878 54139
rect 1066 52485 438878 53051
rect 1066 51397 438878 51963
rect 1066 50309 438878 50875
rect 1066 49221 438878 49787
rect 1066 48133 438878 48699
rect 1066 47045 438878 47611
rect 1066 45957 438878 46523
rect 1066 44869 438878 45435
rect 1066 43781 438878 44347
rect 1066 42693 438878 43259
rect 1066 41605 438878 42171
rect 1066 40517 438878 41083
rect 1066 39429 438878 39995
rect 1066 38341 438878 38907
rect 1066 37253 438878 37819
rect 1066 36165 438878 36731
rect 1066 35077 438878 35643
rect 1066 33989 438878 34555
rect 1066 32901 438878 33467
rect 1066 31813 438878 32379
rect 1066 30725 438878 31291
rect 1066 29637 438878 30203
rect 1066 28549 438878 29115
rect 1066 27461 438878 28027
rect 1066 26373 438878 26939
rect 1066 25285 438878 25851
rect 1066 24197 438878 24763
rect 1066 23109 438878 23675
rect 1066 22021 438878 22587
rect 1066 20933 438878 21499
rect 1066 19845 438878 20411
rect 1066 18757 438878 19323
rect 1066 17669 438878 18235
rect 1066 16581 438878 17147
rect 1066 15493 438878 16059
rect 1066 14405 438878 14971
rect 1066 13317 438878 13883
rect 1066 12229 438878 12795
rect 1066 11141 438878 11707
rect 1066 10053 438878 10619
rect 1066 8965 438878 9531
rect 1066 7877 438878 8443
rect 1066 6789 438878 7355
rect 1066 5701 438878 6267
rect 1066 4613 438878 5179
rect 1066 3525 438878 4091
rect 1066 2437 438878 3003
<< obsli1 >>
rect 1104 2159 438840 557617
<< obsm1 >>
rect 1104 144 439010 557648
<< metal2 >>
rect 6826 559200 6882 560000
rect 10598 559200 10654 560000
rect 14370 559200 14426 560000
rect 18142 559200 18198 560000
rect 21914 559200 21970 560000
rect 25686 559200 25742 560000
rect 29458 559200 29514 560000
rect 33230 559200 33286 560000
rect 37002 559200 37058 560000
rect 40774 559200 40830 560000
rect 44546 559200 44602 560000
rect 48318 559200 48374 560000
rect 52090 559200 52146 560000
rect 55862 559200 55918 560000
rect 59634 559200 59690 560000
rect 63406 559200 63462 560000
rect 67178 559200 67234 560000
rect 70950 559200 71006 560000
rect 74722 559200 74778 560000
rect 78494 559200 78550 560000
rect 82266 559200 82322 560000
rect 86038 559200 86094 560000
rect 89810 559200 89866 560000
rect 93582 559200 93638 560000
rect 97354 559200 97410 560000
rect 101126 559200 101182 560000
rect 104898 559200 104954 560000
rect 108670 559200 108726 560000
rect 112442 559200 112498 560000
rect 116214 559200 116270 560000
rect 119986 559200 120042 560000
rect 123758 559200 123814 560000
rect 127530 559200 127586 560000
rect 131302 559200 131358 560000
rect 135074 559200 135130 560000
rect 138846 559200 138902 560000
rect 142618 559200 142674 560000
rect 146390 559200 146446 560000
rect 150162 559200 150218 560000
rect 153934 559200 153990 560000
rect 157706 559200 157762 560000
rect 161478 559200 161534 560000
rect 165250 559200 165306 560000
rect 169022 559200 169078 560000
rect 172794 559200 172850 560000
rect 176566 559200 176622 560000
rect 180338 559200 180394 560000
rect 184110 559200 184166 560000
rect 187882 559200 187938 560000
rect 191654 559200 191710 560000
rect 195426 559200 195482 560000
rect 199198 559200 199254 560000
rect 202970 559200 203026 560000
rect 206742 559200 206798 560000
rect 210514 559200 210570 560000
rect 214286 559200 214342 560000
rect 218058 559200 218114 560000
rect 221830 559200 221886 560000
rect 225602 559200 225658 560000
rect 229374 559200 229430 560000
rect 233146 559200 233202 560000
rect 236918 559200 236974 560000
rect 240690 559200 240746 560000
rect 244462 559200 244518 560000
rect 248234 559200 248290 560000
rect 252006 559200 252062 560000
rect 255778 559200 255834 560000
rect 259550 559200 259606 560000
rect 263322 559200 263378 560000
rect 267094 559200 267150 560000
rect 270866 559200 270922 560000
rect 274638 559200 274694 560000
rect 278410 559200 278466 560000
rect 282182 559200 282238 560000
rect 285954 559200 286010 560000
rect 289726 559200 289782 560000
rect 293498 559200 293554 560000
rect 297270 559200 297326 560000
rect 301042 559200 301098 560000
rect 304814 559200 304870 560000
rect 308586 559200 308642 560000
rect 312358 559200 312414 560000
rect 316130 559200 316186 560000
rect 319902 559200 319958 560000
rect 323674 559200 323730 560000
rect 327446 559200 327502 560000
rect 331218 559200 331274 560000
rect 334990 559200 335046 560000
rect 338762 559200 338818 560000
rect 342534 559200 342590 560000
rect 346306 559200 346362 560000
rect 350078 559200 350134 560000
rect 353850 559200 353906 560000
rect 357622 559200 357678 560000
rect 361394 559200 361450 560000
rect 365166 559200 365222 560000
rect 368938 559200 368994 560000
rect 372710 559200 372766 560000
rect 376482 559200 376538 560000
rect 380254 559200 380310 560000
rect 384026 559200 384082 560000
rect 387798 559200 387854 560000
rect 391570 559200 391626 560000
rect 395342 559200 395398 560000
rect 399114 559200 399170 560000
rect 402886 559200 402942 560000
rect 406658 559200 406714 560000
rect 410430 559200 410486 560000
rect 414202 559200 414258 560000
rect 417974 559200 418030 560000
rect 421746 559200 421802 560000
rect 425518 559200 425574 560000
rect 429290 559200 429346 560000
rect 433062 559200 433118 560000
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19614 0 19670 800
rect 20442 0 20498 800
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 57702 0 57758 800
rect 58530 0 58586 800
rect 59358 0 59414 800
rect 60186 0 60242 800
rect 61014 0 61070 800
rect 61842 0 61898 800
rect 62670 0 62726 800
rect 63498 0 63554 800
rect 64326 0 64382 800
rect 65154 0 65210 800
rect 65982 0 66038 800
rect 66810 0 66866 800
rect 67638 0 67694 800
rect 68466 0 68522 800
rect 69294 0 69350 800
rect 70122 0 70178 800
rect 70950 0 71006 800
rect 71778 0 71834 800
rect 72606 0 72662 800
rect 73434 0 73490 800
rect 74262 0 74318 800
rect 75090 0 75146 800
rect 75918 0 75974 800
rect 76746 0 76802 800
rect 77574 0 77630 800
rect 78402 0 78458 800
rect 79230 0 79286 800
rect 80058 0 80114 800
rect 80886 0 80942 800
rect 81714 0 81770 800
rect 82542 0 82598 800
rect 83370 0 83426 800
rect 84198 0 84254 800
rect 85026 0 85082 800
rect 85854 0 85910 800
rect 86682 0 86738 800
rect 87510 0 87566 800
rect 88338 0 88394 800
rect 89166 0 89222 800
rect 89994 0 90050 800
rect 90822 0 90878 800
rect 91650 0 91706 800
rect 92478 0 92534 800
rect 93306 0 93362 800
rect 94134 0 94190 800
rect 94962 0 95018 800
rect 95790 0 95846 800
rect 96618 0 96674 800
rect 97446 0 97502 800
rect 98274 0 98330 800
rect 99102 0 99158 800
rect 99930 0 99986 800
rect 100758 0 100814 800
rect 101586 0 101642 800
rect 102414 0 102470 800
rect 103242 0 103298 800
rect 104070 0 104126 800
rect 104898 0 104954 800
rect 105726 0 105782 800
rect 106554 0 106610 800
rect 107382 0 107438 800
rect 108210 0 108266 800
rect 109038 0 109094 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113178 0 113234 800
rect 114006 0 114062 800
rect 114834 0 114890 800
rect 115662 0 115718 800
rect 116490 0 116546 800
rect 117318 0 117374 800
rect 118146 0 118202 800
rect 118974 0 119030 800
rect 119802 0 119858 800
rect 120630 0 120686 800
rect 121458 0 121514 800
rect 122286 0 122342 800
rect 123114 0 123170 800
rect 123942 0 123998 800
rect 124770 0 124826 800
rect 125598 0 125654 800
rect 126426 0 126482 800
rect 127254 0 127310 800
rect 128082 0 128138 800
rect 128910 0 128966 800
rect 129738 0 129794 800
rect 130566 0 130622 800
rect 131394 0 131450 800
rect 132222 0 132278 800
rect 133050 0 133106 800
rect 133878 0 133934 800
rect 134706 0 134762 800
rect 135534 0 135590 800
rect 136362 0 136418 800
rect 137190 0 137246 800
rect 138018 0 138074 800
rect 138846 0 138902 800
rect 139674 0 139730 800
rect 140502 0 140558 800
rect 141330 0 141386 800
rect 142158 0 142214 800
rect 142986 0 143042 800
rect 143814 0 143870 800
rect 144642 0 144698 800
rect 145470 0 145526 800
rect 146298 0 146354 800
rect 147126 0 147182 800
rect 147954 0 148010 800
rect 148782 0 148838 800
rect 149610 0 149666 800
rect 150438 0 150494 800
rect 151266 0 151322 800
rect 152094 0 152150 800
rect 152922 0 152978 800
rect 153750 0 153806 800
rect 154578 0 154634 800
rect 155406 0 155462 800
rect 156234 0 156290 800
rect 157062 0 157118 800
rect 157890 0 157946 800
rect 158718 0 158774 800
rect 159546 0 159602 800
rect 160374 0 160430 800
rect 161202 0 161258 800
rect 162030 0 162086 800
rect 162858 0 162914 800
rect 163686 0 163742 800
rect 164514 0 164570 800
rect 165342 0 165398 800
rect 166170 0 166226 800
rect 166998 0 167054 800
rect 167826 0 167882 800
rect 168654 0 168710 800
rect 169482 0 169538 800
rect 170310 0 170366 800
rect 171138 0 171194 800
rect 171966 0 172022 800
rect 172794 0 172850 800
rect 173622 0 173678 800
rect 174450 0 174506 800
rect 175278 0 175334 800
rect 176106 0 176162 800
rect 176934 0 176990 800
rect 177762 0 177818 800
rect 178590 0 178646 800
rect 179418 0 179474 800
rect 180246 0 180302 800
rect 181074 0 181130 800
rect 181902 0 181958 800
rect 182730 0 182786 800
rect 183558 0 183614 800
rect 184386 0 184442 800
rect 185214 0 185270 800
rect 186042 0 186098 800
rect 186870 0 186926 800
rect 187698 0 187754 800
rect 188526 0 188582 800
rect 189354 0 189410 800
rect 190182 0 190238 800
rect 191010 0 191066 800
rect 191838 0 191894 800
rect 192666 0 192722 800
rect 193494 0 193550 800
rect 194322 0 194378 800
rect 195150 0 195206 800
rect 195978 0 196034 800
rect 196806 0 196862 800
rect 197634 0 197690 800
rect 198462 0 198518 800
rect 199290 0 199346 800
rect 200118 0 200174 800
rect 200946 0 201002 800
rect 201774 0 201830 800
rect 202602 0 202658 800
rect 203430 0 203486 800
rect 204258 0 204314 800
rect 205086 0 205142 800
rect 205914 0 205970 800
rect 206742 0 206798 800
rect 207570 0 207626 800
rect 208398 0 208454 800
rect 209226 0 209282 800
rect 210054 0 210110 800
rect 210882 0 210938 800
rect 211710 0 211766 800
rect 212538 0 212594 800
rect 213366 0 213422 800
rect 214194 0 214250 800
rect 215022 0 215078 800
rect 215850 0 215906 800
rect 216678 0 216734 800
rect 217506 0 217562 800
rect 218334 0 218390 800
rect 219162 0 219218 800
rect 219990 0 220046 800
rect 220818 0 220874 800
rect 221646 0 221702 800
rect 222474 0 222530 800
rect 223302 0 223358 800
rect 224130 0 224186 800
rect 224958 0 225014 800
rect 225786 0 225842 800
rect 226614 0 226670 800
rect 227442 0 227498 800
rect 228270 0 228326 800
rect 229098 0 229154 800
rect 229926 0 229982 800
rect 230754 0 230810 800
rect 231582 0 231638 800
rect 232410 0 232466 800
rect 233238 0 233294 800
rect 234066 0 234122 800
rect 234894 0 234950 800
rect 235722 0 235778 800
rect 236550 0 236606 800
rect 237378 0 237434 800
rect 238206 0 238262 800
rect 239034 0 239090 800
rect 239862 0 239918 800
rect 240690 0 240746 800
rect 241518 0 241574 800
rect 242346 0 242402 800
rect 243174 0 243230 800
rect 244002 0 244058 800
rect 244830 0 244886 800
rect 245658 0 245714 800
rect 246486 0 246542 800
rect 247314 0 247370 800
rect 248142 0 248198 800
rect 248970 0 249026 800
rect 249798 0 249854 800
rect 250626 0 250682 800
rect 251454 0 251510 800
rect 252282 0 252338 800
rect 253110 0 253166 800
rect 253938 0 253994 800
rect 254766 0 254822 800
rect 255594 0 255650 800
rect 256422 0 256478 800
rect 257250 0 257306 800
rect 258078 0 258134 800
rect 258906 0 258962 800
rect 259734 0 259790 800
rect 260562 0 260618 800
rect 261390 0 261446 800
rect 262218 0 262274 800
rect 263046 0 263102 800
rect 263874 0 263930 800
rect 264702 0 264758 800
rect 265530 0 265586 800
rect 266358 0 266414 800
rect 267186 0 267242 800
rect 268014 0 268070 800
rect 268842 0 268898 800
rect 269670 0 269726 800
rect 270498 0 270554 800
rect 271326 0 271382 800
rect 272154 0 272210 800
rect 272982 0 273038 800
rect 273810 0 273866 800
rect 274638 0 274694 800
rect 275466 0 275522 800
rect 276294 0 276350 800
rect 277122 0 277178 800
rect 277950 0 278006 800
rect 278778 0 278834 800
rect 279606 0 279662 800
rect 280434 0 280490 800
rect 281262 0 281318 800
rect 282090 0 282146 800
rect 282918 0 282974 800
rect 283746 0 283802 800
rect 284574 0 284630 800
rect 285402 0 285458 800
rect 286230 0 286286 800
rect 287058 0 287114 800
rect 287886 0 287942 800
rect 288714 0 288770 800
rect 289542 0 289598 800
rect 290370 0 290426 800
rect 291198 0 291254 800
rect 292026 0 292082 800
rect 292854 0 292910 800
rect 293682 0 293738 800
rect 294510 0 294566 800
rect 295338 0 295394 800
rect 296166 0 296222 800
rect 296994 0 297050 800
rect 297822 0 297878 800
rect 298650 0 298706 800
rect 299478 0 299534 800
rect 300306 0 300362 800
rect 301134 0 301190 800
rect 301962 0 302018 800
rect 302790 0 302846 800
rect 303618 0 303674 800
rect 304446 0 304502 800
rect 305274 0 305330 800
rect 306102 0 306158 800
rect 306930 0 306986 800
rect 307758 0 307814 800
rect 308586 0 308642 800
rect 309414 0 309470 800
rect 310242 0 310298 800
rect 311070 0 311126 800
rect 311898 0 311954 800
rect 312726 0 312782 800
rect 313554 0 313610 800
rect 314382 0 314438 800
rect 315210 0 315266 800
rect 316038 0 316094 800
rect 316866 0 316922 800
rect 317694 0 317750 800
rect 318522 0 318578 800
rect 319350 0 319406 800
rect 320178 0 320234 800
rect 321006 0 321062 800
rect 321834 0 321890 800
rect 322662 0 322718 800
rect 323490 0 323546 800
rect 324318 0 324374 800
rect 325146 0 325202 800
rect 325974 0 326030 800
rect 326802 0 326858 800
rect 327630 0 327686 800
rect 328458 0 328514 800
rect 329286 0 329342 800
rect 330114 0 330170 800
rect 330942 0 330998 800
rect 331770 0 331826 800
rect 332598 0 332654 800
rect 333426 0 333482 800
rect 334254 0 334310 800
rect 335082 0 335138 800
rect 335910 0 335966 800
rect 336738 0 336794 800
rect 337566 0 337622 800
rect 338394 0 338450 800
rect 339222 0 339278 800
rect 340050 0 340106 800
rect 340878 0 340934 800
rect 341706 0 341762 800
rect 342534 0 342590 800
rect 343362 0 343418 800
rect 344190 0 344246 800
rect 345018 0 345074 800
rect 345846 0 345902 800
rect 346674 0 346730 800
rect 347502 0 347558 800
rect 348330 0 348386 800
rect 349158 0 349214 800
rect 349986 0 350042 800
rect 350814 0 350870 800
rect 351642 0 351698 800
rect 352470 0 352526 800
rect 353298 0 353354 800
rect 354126 0 354182 800
rect 354954 0 355010 800
rect 355782 0 355838 800
rect 356610 0 356666 800
rect 357438 0 357494 800
rect 358266 0 358322 800
rect 359094 0 359150 800
rect 359922 0 359978 800
rect 360750 0 360806 800
rect 361578 0 361634 800
rect 362406 0 362462 800
rect 363234 0 363290 800
rect 364062 0 364118 800
rect 364890 0 364946 800
rect 365718 0 365774 800
rect 366546 0 366602 800
rect 367374 0 367430 800
rect 368202 0 368258 800
rect 369030 0 369086 800
rect 369858 0 369914 800
rect 370686 0 370742 800
rect 371514 0 371570 800
rect 372342 0 372398 800
rect 373170 0 373226 800
rect 373998 0 374054 800
rect 374826 0 374882 800
rect 375654 0 375710 800
rect 376482 0 376538 800
rect 377310 0 377366 800
rect 378138 0 378194 800
rect 378966 0 379022 800
rect 379794 0 379850 800
rect 380622 0 380678 800
rect 381450 0 381506 800
rect 382278 0 382334 800
rect 383106 0 383162 800
rect 383934 0 383990 800
rect 384762 0 384818 800
rect 385590 0 385646 800
rect 386418 0 386474 800
rect 387246 0 387302 800
rect 388074 0 388130 800
rect 388902 0 388958 800
rect 389730 0 389786 800
rect 390558 0 390614 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394698 0 394754 800
rect 395526 0 395582 800
rect 396354 0 396410 800
rect 397182 0 397238 800
rect 398010 0 398066 800
rect 398838 0 398894 800
rect 399666 0 399722 800
rect 400494 0 400550 800
rect 401322 0 401378 800
rect 402150 0 402206 800
rect 402978 0 403034 800
rect 403806 0 403862 800
rect 404634 0 404690 800
rect 405462 0 405518 800
rect 406290 0 406346 800
rect 407118 0 407174 800
rect 407946 0 408002 800
rect 408774 0 408830 800
rect 409602 0 409658 800
rect 410430 0 410486 800
rect 411258 0 411314 800
rect 412086 0 412142 800
rect 412914 0 412970 800
rect 413742 0 413798 800
rect 414570 0 414626 800
rect 415398 0 415454 800
rect 416226 0 416282 800
rect 417054 0 417110 800
rect 417882 0 417938 800
rect 418710 0 418766 800
rect 419538 0 419594 800
rect 420366 0 420422 800
rect 421194 0 421250 800
rect 422022 0 422078 800
rect 422850 0 422906 800
rect 423678 0 423734 800
<< obsm2 >>
rect 1400 559144 6770 559314
rect 6938 559144 10542 559314
rect 10710 559144 14314 559314
rect 14482 559144 18086 559314
rect 18254 559144 21858 559314
rect 22026 559144 25630 559314
rect 25798 559144 29402 559314
rect 29570 559144 33174 559314
rect 33342 559144 36946 559314
rect 37114 559144 40718 559314
rect 40886 559144 44490 559314
rect 44658 559144 48262 559314
rect 48430 559144 52034 559314
rect 52202 559144 55806 559314
rect 55974 559144 59578 559314
rect 59746 559144 63350 559314
rect 63518 559144 67122 559314
rect 67290 559144 70894 559314
rect 71062 559144 74666 559314
rect 74834 559144 78438 559314
rect 78606 559144 82210 559314
rect 82378 559144 85982 559314
rect 86150 559144 89754 559314
rect 89922 559144 93526 559314
rect 93694 559144 97298 559314
rect 97466 559144 101070 559314
rect 101238 559144 104842 559314
rect 105010 559144 108614 559314
rect 108782 559144 112386 559314
rect 112554 559144 116158 559314
rect 116326 559144 119930 559314
rect 120098 559144 123702 559314
rect 123870 559144 127474 559314
rect 127642 559144 131246 559314
rect 131414 559144 135018 559314
rect 135186 559144 138790 559314
rect 138958 559144 142562 559314
rect 142730 559144 146334 559314
rect 146502 559144 150106 559314
rect 150274 559144 153878 559314
rect 154046 559144 157650 559314
rect 157818 559144 161422 559314
rect 161590 559144 165194 559314
rect 165362 559144 168966 559314
rect 169134 559144 172738 559314
rect 172906 559144 176510 559314
rect 176678 559144 180282 559314
rect 180450 559144 184054 559314
rect 184222 559144 187826 559314
rect 187994 559144 191598 559314
rect 191766 559144 195370 559314
rect 195538 559144 199142 559314
rect 199310 559144 202914 559314
rect 203082 559144 206686 559314
rect 206854 559144 210458 559314
rect 210626 559144 214230 559314
rect 214398 559144 218002 559314
rect 218170 559144 221774 559314
rect 221942 559144 225546 559314
rect 225714 559144 229318 559314
rect 229486 559144 233090 559314
rect 233258 559144 236862 559314
rect 237030 559144 240634 559314
rect 240802 559144 244406 559314
rect 244574 559144 248178 559314
rect 248346 559144 251950 559314
rect 252118 559144 255722 559314
rect 255890 559144 259494 559314
rect 259662 559144 263266 559314
rect 263434 559144 267038 559314
rect 267206 559144 270810 559314
rect 270978 559144 274582 559314
rect 274750 559144 278354 559314
rect 278522 559144 282126 559314
rect 282294 559144 285898 559314
rect 286066 559144 289670 559314
rect 289838 559144 293442 559314
rect 293610 559144 297214 559314
rect 297382 559144 300986 559314
rect 301154 559144 304758 559314
rect 304926 559144 308530 559314
rect 308698 559144 312302 559314
rect 312470 559144 316074 559314
rect 316242 559144 319846 559314
rect 320014 559144 323618 559314
rect 323786 559144 327390 559314
rect 327558 559144 331162 559314
rect 331330 559144 334934 559314
rect 335102 559144 338706 559314
rect 338874 559144 342478 559314
rect 342646 559144 346250 559314
rect 346418 559144 350022 559314
rect 350190 559144 353794 559314
rect 353962 559144 357566 559314
rect 357734 559144 361338 559314
rect 361506 559144 365110 559314
rect 365278 559144 368882 559314
rect 369050 559144 372654 559314
rect 372822 559144 376426 559314
rect 376594 559144 380198 559314
rect 380366 559144 383970 559314
rect 384138 559144 387742 559314
rect 387910 559144 391514 559314
rect 391682 559144 395286 559314
rect 395454 559144 399058 559314
rect 399226 559144 402830 559314
rect 402998 559144 406602 559314
rect 406770 559144 410374 559314
rect 410542 559144 414146 559314
rect 414314 559144 417918 559314
rect 418086 559144 421690 559314
rect 421858 559144 425462 559314
rect 425630 559144 429234 559314
rect 429402 559144 433006 559314
rect 433174 559144 439006 559314
rect 1400 856 439006 559144
rect 1400 138 16246 856
rect 16414 138 17074 856
rect 17242 138 17902 856
rect 18070 138 18730 856
rect 18898 138 19558 856
rect 19726 138 20386 856
rect 20554 138 21214 856
rect 21382 138 22042 856
rect 22210 138 22870 856
rect 23038 138 23698 856
rect 23866 138 24526 856
rect 24694 138 25354 856
rect 25522 138 26182 856
rect 26350 138 27010 856
rect 27178 138 27838 856
rect 28006 138 28666 856
rect 28834 138 29494 856
rect 29662 138 30322 856
rect 30490 138 31150 856
rect 31318 138 31978 856
rect 32146 138 32806 856
rect 32974 138 33634 856
rect 33802 138 34462 856
rect 34630 138 35290 856
rect 35458 138 36118 856
rect 36286 138 36946 856
rect 37114 138 37774 856
rect 37942 138 38602 856
rect 38770 138 39430 856
rect 39598 138 40258 856
rect 40426 138 41086 856
rect 41254 138 41914 856
rect 42082 138 42742 856
rect 42910 138 43570 856
rect 43738 138 44398 856
rect 44566 138 45226 856
rect 45394 138 46054 856
rect 46222 138 46882 856
rect 47050 138 47710 856
rect 47878 138 48538 856
rect 48706 138 49366 856
rect 49534 138 50194 856
rect 50362 138 51022 856
rect 51190 138 51850 856
rect 52018 138 52678 856
rect 52846 138 53506 856
rect 53674 138 54334 856
rect 54502 138 55162 856
rect 55330 138 55990 856
rect 56158 138 56818 856
rect 56986 138 57646 856
rect 57814 138 58474 856
rect 58642 138 59302 856
rect 59470 138 60130 856
rect 60298 138 60958 856
rect 61126 138 61786 856
rect 61954 138 62614 856
rect 62782 138 63442 856
rect 63610 138 64270 856
rect 64438 138 65098 856
rect 65266 138 65926 856
rect 66094 138 66754 856
rect 66922 138 67582 856
rect 67750 138 68410 856
rect 68578 138 69238 856
rect 69406 138 70066 856
rect 70234 138 70894 856
rect 71062 138 71722 856
rect 71890 138 72550 856
rect 72718 138 73378 856
rect 73546 138 74206 856
rect 74374 138 75034 856
rect 75202 138 75862 856
rect 76030 138 76690 856
rect 76858 138 77518 856
rect 77686 138 78346 856
rect 78514 138 79174 856
rect 79342 138 80002 856
rect 80170 138 80830 856
rect 80998 138 81658 856
rect 81826 138 82486 856
rect 82654 138 83314 856
rect 83482 138 84142 856
rect 84310 138 84970 856
rect 85138 138 85798 856
rect 85966 138 86626 856
rect 86794 138 87454 856
rect 87622 138 88282 856
rect 88450 138 89110 856
rect 89278 138 89938 856
rect 90106 138 90766 856
rect 90934 138 91594 856
rect 91762 138 92422 856
rect 92590 138 93250 856
rect 93418 138 94078 856
rect 94246 138 94906 856
rect 95074 138 95734 856
rect 95902 138 96562 856
rect 96730 138 97390 856
rect 97558 138 98218 856
rect 98386 138 99046 856
rect 99214 138 99874 856
rect 100042 138 100702 856
rect 100870 138 101530 856
rect 101698 138 102358 856
rect 102526 138 103186 856
rect 103354 138 104014 856
rect 104182 138 104842 856
rect 105010 138 105670 856
rect 105838 138 106498 856
rect 106666 138 107326 856
rect 107494 138 108154 856
rect 108322 138 108982 856
rect 109150 138 109810 856
rect 109978 138 110638 856
rect 110806 138 111466 856
rect 111634 138 112294 856
rect 112462 138 113122 856
rect 113290 138 113950 856
rect 114118 138 114778 856
rect 114946 138 115606 856
rect 115774 138 116434 856
rect 116602 138 117262 856
rect 117430 138 118090 856
rect 118258 138 118918 856
rect 119086 138 119746 856
rect 119914 138 120574 856
rect 120742 138 121402 856
rect 121570 138 122230 856
rect 122398 138 123058 856
rect 123226 138 123886 856
rect 124054 138 124714 856
rect 124882 138 125542 856
rect 125710 138 126370 856
rect 126538 138 127198 856
rect 127366 138 128026 856
rect 128194 138 128854 856
rect 129022 138 129682 856
rect 129850 138 130510 856
rect 130678 138 131338 856
rect 131506 138 132166 856
rect 132334 138 132994 856
rect 133162 138 133822 856
rect 133990 138 134650 856
rect 134818 138 135478 856
rect 135646 138 136306 856
rect 136474 138 137134 856
rect 137302 138 137962 856
rect 138130 138 138790 856
rect 138958 138 139618 856
rect 139786 138 140446 856
rect 140614 138 141274 856
rect 141442 138 142102 856
rect 142270 138 142930 856
rect 143098 138 143758 856
rect 143926 138 144586 856
rect 144754 138 145414 856
rect 145582 138 146242 856
rect 146410 138 147070 856
rect 147238 138 147898 856
rect 148066 138 148726 856
rect 148894 138 149554 856
rect 149722 138 150382 856
rect 150550 138 151210 856
rect 151378 138 152038 856
rect 152206 138 152866 856
rect 153034 138 153694 856
rect 153862 138 154522 856
rect 154690 138 155350 856
rect 155518 138 156178 856
rect 156346 138 157006 856
rect 157174 138 157834 856
rect 158002 138 158662 856
rect 158830 138 159490 856
rect 159658 138 160318 856
rect 160486 138 161146 856
rect 161314 138 161974 856
rect 162142 138 162802 856
rect 162970 138 163630 856
rect 163798 138 164458 856
rect 164626 138 165286 856
rect 165454 138 166114 856
rect 166282 138 166942 856
rect 167110 138 167770 856
rect 167938 138 168598 856
rect 168766 138 169426 856
rect 169594 138 170254 856
rect 170422 138 171082 856
rect 171250 138 171910 856
rect 172078 138 172738 856
rect 172906 138 173566 856
rect 173734 138 174394 856
rect 174562 138 175222 856
rect 175390 138 176050 856
rect 176218 138 176878 856
rect 177046 138 177706 856
rect 177874 138 178534 856
rect 178702 138 179362 856
rect 179530 138 180190 856
rect 180358 138 181018 856
rect 181186 138 181846 856
rect 182014 138 182674 856
rect 182842 138 183502 856
rect 183670 138 184330 856
rect 184498 138 185158 856
rect 185326 138 185986 856
rect 186154 138 186814 856
rect 186982 138 187642 856
rect 187810 138 188470 856
rect 188638 138 189298 856
rect 189466 138 190126 856
rect 190294 138 190954 856
rect 191122 138 191782 856
rect 191950 138 192610 856
rect 192778 138 193438 856
rect 193606 138 194266 856
rect 194434 138 195094 856
rect 195262 138 195922 856
rect 196090 138 196750 856
rect 196918 138 197578 856
rect 197746 138 198406 856
rect 198574 138 199234 856
rect 199402 138 200062 856
rect 200230 138 200890 856
rect 201058 138 201718 856
rect 201886 138 202546 856
rect 202714 138 203374 856
rect 203542 138 204202 856
rect 204370 138 205030 856
rect 205198 138 205858 856
rect 206026 138 206686 856
rect 206854 138 207514 856
rect 207682 138 208342 856
rect 208510 138 209170 856
rect 209338 138 209998 856
rect 210166 138 210826 856
rect 210994 138 211654 856
rect 211822 138 212482 856
rect 212650 138 213310 856
rect 213478 138 214138 856
rect 214306 138 214966 856
rect 215134 138 215794 856
rect 215962 138 216622 856
rect 216790 138 217450 856
rect 217618 138 218278 856
rect 218446 138 219106 856
rect 219274 138 219934 856
rect 220102 138 220762 856
rect 220930 138 221590 856
rect 221758 138 222418 856
rect 222586 138 223246 856
rect 223414 138 224074 856
rect 224242 138 224902 856
rect 225070 138 225730 856
rect 225898 138 226558 856
rect 226726 138 227386 856
rect 227554 138 228214 856
rect 228382 138 229042 856
rect 229210 138 229870 856
rect 230038 138 230698 856
rect 230866 138 231526 856
rect 231694 138 232354 856
rect 232522 138 233182 856
rect 233350 138 234010 856
rect 234178 138 234838 856
rect 235006 138 235666 856
rect 235834 138 236494 856
rect 236662 138 237322 856
rect 237490 138 238150 856
rect 238318 138 238978 856
rect 239146 138 239806 856
rect 239974 138 240634 856
rect 240802 138 241462 856
rect 241630 138 242290 856
rect 242458 138 243118 856
rect 243286 138 243946 856
rect 244114 138 244774 856
rect 244942 138 245602 856
rect 245770 138 246430 856
rect 246598 138 247258 856
rect 247426 138 248086 856
rect 248254 138 248914 856
rect 249082 138 249742 856
rect 249910 138 250570 856
rect 250738 138 251398 856
rect 251566 138 252226 856
rect 252394 138 253054 856
rect 253222 138 253882 856
rect 254050 138 254710 856
rect 254878 138 255538 856
rect 255706 138 256366 856
rect 256534 138 257194 856
rect 257362 138 258022 856
rect 258190 138 258850 856
rect 259018 138 259678 856
rect 259846 138 260506 856
rect 260674 138 261334 856
rect 261502 138 262162 856
rect 262330 138 262990 856
rect 263158 138 263818 856
rect 263986 138 264646 856
rect 264814 138 265474 856
rect 265642 138 266302 856
rect 266470 138 267130 856
rect 267298 138 267958 856
rect 268126 138 268786 856
rect 268954 138 269614 856
rect 269782 138 270442 856
rect 270610 138 271270 856
rect 271438 138 272098 856
rect 272266 138 272926 856
rect 273094 138 273754 856
rect 273922 138 274582 856
rect 274750 138 275410 856
rect 275578 138 276238 856
rect 276406 138 277066 856
rect 277234 138 277894 856
rect 278062 138 278722 856
rect 278890 138 279550 856
rect 279718 138 280378 856
rect 280546 138 281206 856
rect 281374 138 282034 856
rect 282202 138 282862 856
rect 283030 138 283690 856
rect 283858 138 284518 856
rect 284686 138 285346 856
rect 285514 138 286174 856
rect 286342 138 287002 856
rect 287170 138 287830 856
rect 287998 138 288658 856
rect 288826 138 289486 856
rect 289654 138 290314 856
rect 290482 138 291142 856
rect 291310 138 291970 856
rect 292138 138 292798 856
rect 292966 138 293626 856
rect 293794 138 294454 856
rect 294622 138 295282 856
rect 295450 138 296110 856
rect 296278 138 296938 856
rect 297106 138 297766 856
rect 297934 138 298594 856
rect 298762 138 299422 856
rect 299590 138 300250 856
rect 300418 138 301078 856
rect 301246 138 301906 856
rect 302074 138 302734 856
rect 302902 138 303562 856
rect 303730 138 304390 856
rect 304558 138 305218 856
rect 305386 138 306046 856
rect 306214 138 306874 856
rect 307042 138 307702 856
rect 307870 138 308530 856
rect 308698 138 309358 856
rect 309526 138 310186 856
rect 310354 138 311014 856
rect 311182 138 311842 856
rect 312010 138 312670 856
rect 312838 138 313498 856
rect 313666 138 314326 856
rect 314494 138 315154 856
rect 315322 138 315982 856
rect 316150 138 316810 856
rect 316978 138 317638 856
rect 317806 138 318466 856
rect 318634 138 319294 856
rect 319462 138 320122 856
rect 320290 138 320950 856
rect 321118 138 321778 856
rect 321946 138 322606 856
rect 322774 138 323434 856
rect 323602 138 324262 856
rect 324430 138 325090 856
rect 325258 138 325918 856
rect 326086 138 326746 856
rect 326914 138 327574 856
rect 327742 138 328402 856
rect 328570 138 329230 856
rect 329398 138 330058 856
rect 330226 138 330886 856
rect 331054 138 331714 856
rect 331882 138 332542 856
rect 332710 138 333370 856
rect 333538 138 334198 856
rect 334366 138 335026 856
rect 335194 138 335854 856
rect 336022 138 336682 856
rect 336850 138 337510 856
rect 337678 138 338338 856
rect 338506 138 339166 856
rect 339334 138 339994 856
rect 340162 138 340822 856
rect 340990 138 341650 856
rect 341818 138 342478 856
rect 342646 138 343306 856
rect 343474 138 344134 856
rect 344302 138 344962 856
rect 345130 138 345790 856
rect 345958 138 346618 856
rect 346786 138 347446 856
rect 347614 138 348274 856
rect 348442 138 349102 856
rect 349270 138 349930 856
rect 350098 138 350758 856
rect 350926 138 351586 856
rect 351754 138 352414 856
rect 352582 138 353242 856
rect 353410 138 354070 856
rect 354238 138 354898 856
rect 355066 138 355726 856
rect 355894 138 356554 856
rect 356722 138 357382 856
rect 357550 138 358210 856
rect 358378 138 359038 856
rect 359206 138 359866 856
rect 360034 138 360694 856
rect 360862 138 361522 856
rect 361690 138 362350 856
rect 362518 138 363178 856
rect 363346 138 364006 856
rect 364174 138 364834 856
rect 365002 138 365662 856
rect 365830 138 366490 856
rect 366658 138 367318 856
rect 367486 138 368146 856
rect 368314 138 368974 856
rect 369142 138 369802 856
rect 369970 138 370630 856
rect 370798 138 371458 856
rect 371626 138 372286 856
rect 372454 138 373114 856
rect 373282 138 373942 856
rect 374110 138 374770 856
rect 374938 138 375598 856
rect 375766 138 376426 856
rect 376594 138 377254 856
rect 377422 138 378082 856
rect 378250 138 378910 856
rect 379078 138 379738 856
rect 379906 138 380566 856
rect 380734 138 381394 856
rect 381562 138 382222 856
rect 382390 138 383050 856
rect 383218 138 383878 856
rect 384046 138 384706 856
rect 384874 138 385534 856
rect 385702 138 386362 856
rect 386530 138 387190 856
rect 387358 138 388018 856
rect 388186 138 388846 856
rect 389014 138 389674 856
rect 389842 138 390502 856
rect 390670 138 391330 856
rect 391498 138 392158 856
rect 392326 138 392986 856
rect 393154 138 393814 856
rect 393982 138 394642 856
rect 394810 138 395470 856
rect 395638 138 396298 856
rect 396466 138 397126 856
rect 397294 138 397954 856
rect 398122 138 398782 856
rect 398950 138 399610 856
rect 399778 138 400438 856
rect 400606 138 401266 856
rect 401434 138 402094 856
rect 402262 138 402922 856
rect 403090 138 403750 856
rect 403918 138 404578 856
rect 404746 138 405406 856
rect 405574 138 406234 856
rect 406402 138 407062 856
rect 407230 138 407890 856
rect 408058 138 408718 856
rect 408886 138 409546 856
rect 409714 138 410374 856
rect 410542 138 411202 856
rect 411370 138 412030 856
rect 412198 138 412858 856
rect 413026 138 413686 856
rect 413854 138 414514 856
rect 414682 138 415342 856
rect 415510 138 416170 856
rect 416338 138 416998 856
rect 417166 138 417826 856
rect 417994 138 418654 856
rect 418822 138 419482 856
rect 419650 138 420310 856
rect 420478 138 421138 856
rect 421306 138 421966 856
rect 422134 138 422794 856
rect 422962 138 423622 856
rect 423790 138 439006 856
<< obsm3 >>
rect 2865 443 439011 557633
<< metal4 >>
rect 4208 2128 4528 557648
rect 19568 2128 19888 557648
rect 34928 2128 35248 557648
rect 50288 2128 50608 557648
rect 65648 2128 65968 557648
rect 81008 2128 81328 557648
rect 96368 2128 96688 557648
rect 111728 2128 112048 557648
rect 127088 2128 127408 557648
rect 142448 2128 142768 557648
rect 157808 2128 158128 557648
rect 173168 2128 173488 557648
rect 188528 2128 188848 557648
rect 203888 2128 204208 557648
rect 219248 2128 219568 557648
rect 234608 2128 234928 557648
rect 249968 2128 250288 557648
rect 265328 2128 265648 557648
rect 280688 2128 281008 557648
rect 296048 2128 296368 557648
rect 311408 2128 311728 557648
rect 326768 2128 327088 557648
rect 342128 2128 342448 557648
rect 357488 2128 357808 557648
rect 372848 2128 373168 557648
rect 388208 2128 388528 557648
rect 403568 2128 403888 557648
rect 418928 2128 419248 557648
rect 434288 2128 434608 557648
<< obsm4 >>
rect 3003 2048 4128 552397
rect 4608 2048 19488 552397
rect 19968 2048 34848 552397
rect 35328 2048 50208 552397
rect 50688 2048 65568 552397
rect 66048 2048 80928 552397
rect 81408 2048 96288 552397
rect 96768 2048 111648 552397
rect 112128 2048 127008 552397
rect 127488 2048 142368 552397
rect 142848 2048 157728 552397
rect 158208 2048 173088 552397
rect 173568 2048 188448 552397
rect 188928 2048 203808 552397
rect 204288 2048 219168 552397
rect 219648 2048 234528 552397
rect 235008 2048 249888 552397
rect 250368 2048 265248 552397
rect 265728 2048 280608 552397
rect 281088 2048 295968 552397
rect 296448 2048 311328 552397
rect 311808 2048 326688 552397
rect 327168 2048 342048 552397
rect 342528 2048 357408 552397
rect 357888 2048 372768 552397
rect 373248 2048 388128 552397
rect 388608 2048 403488 552397
rect 403968 2048 418848 552397
rect 419328 2048 434208 552397
rect 434688 2048 436205 552397
rect 3003 443 436205 2048
<< labels >>
rlabel metal2 s 6826 559200 6882 560000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 119986 559200 120042 560000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 131302 559200 131358 560000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 142618 559200 142674 560000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 153934 559200 153990 560000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 165250 559200 165306 560000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 176566 559200 176622 560000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 187882 559200 187938 560000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 199198 559200 199254 560000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 210514 559200 210570 560000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 221830 559200 221886 560000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 18142 559200 18198 560000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 233146 559200 233202 560000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 244462 559200 244518 560000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 255778 559200 255834 560000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 267094 559200 267150 560000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 278410 559200 278466 560000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 289726 559200 289782 560000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 301042 559200 301098 560000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 312358 559200 312414 560000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 323674 559200 323730 560000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 334990 559200 335046 560000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 29458 559200 29514 560000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 346306 559200 346362 560000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 357622 559200 357678 560000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 368938 559200 368994 560000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 380254 559200 380310 560000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 391570 559200 391626 560000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 402886 559200 402942 560000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 414202 559200 414258 560000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 425518 559200 425574 560000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 40774 559200 40830 560000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 52090 559200 52146 560000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 63406 559200 63462 560000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 74722 559200 74778 560000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 86038 559200 86094 560000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 97354 559200 97410 560000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 108670 559200 108726 560000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 10598 559200 10654 560000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 123758 559200 123814 560000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 135074 559200 135130 560000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 146390 559200 146446 560000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 157706 559200 157762 560000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 169022 559200 169078 560000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 180338 559200 180394 560000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 191654 559200 191710 560000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 202970 559200 203026 560000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 214286 559200 214342 560000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 225602 559200 225658 560000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 21914 559200 21970 560000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 236918 559200 236974 560000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 248234 559200 248290 560000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 259550 559200 259606 560000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 270866 559200 270922 560000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 282182 559200 282238 560000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 293498 559200 293554 560000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 304814 559200 304870 560000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 316130 559200 316186 560000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 327446 559200 327502 560000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 338762 559200 338818 560000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 33230 559200 33286 560000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 350078 559200 350134 560000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 361394 559200 361450 560000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 372710 559200 372766 560000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 384026 559200 384082 560000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 395342 559200 395398 560000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 406658 559200 406714 560000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 417974 559200 418030 560000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 429290 559200 429346 560000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 44546 559200 44602 560000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 55862 559200 55918 560000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 67178 559200 67234 560000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 78494 559200 78550 560000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 89810 559200 89866 560000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 101126 559200 101182 560000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 112442 559200 112498 560000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 14370 559200 14426 560000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 127530 559200 127586 560000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 138846 559200 138902 560000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 150162 559200 150218 560000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 161478 559200 161534 560000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 172794 559200 172850 560000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 184110 559200 184166 560000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 195426 559200 195482 560000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 206742 559200 206798 560000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 218058 559200 218114 560000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 229374 559200 229430 560000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 25686 559200 25742 560000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 240690 559200 240746 560000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 252006 559200 252062 560000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 263322 559200 263378 560000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 274638 559200 274694 560000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 285954 559200 286010 560000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 297270 559200 297326 560000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 308586 559200 308642 560000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 319902 559200 319958 560000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 331218 559200 331274 560000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 342534 559200 342590 560000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 37002 559200 37058 560000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 353850 559200 353906 560000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 365166 559200 365222 560000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 376482 559200 376538 560000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 387798 559200 387854 560000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 399114 559200 399170 560000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 410430 559200 410486 560000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 421746 559200 421802 560000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 433062 559200 433118 560000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 48318 559200 48374 560000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 59634 559200 59690 560000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 70950 559200 71006 560000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 82266 559200 82322 560000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 93582 559200 93638 560000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 104898 559200 104954 560000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 116214 559200 116270 560000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 422022 0 422078 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 422850 0 422906 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 423678 0 423734 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 352470 0 352526 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 359922 0 359978 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 362406 0 362462 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 364890 0 364946 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 367374 0 367430 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 369858 0 369914 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 374826 0 374882 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 377310 0 377366 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 379794 0 379850 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 382278 0 382334 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 384762 0 384818 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 387246 0 387302 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 389730 0 389786 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 397182 0 397238 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 399666 0 399722 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 402150 0 402206 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 404634 0 404690 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 407118 0 407174 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 409602 0 409658 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 412086 0 412142 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 414570 0 414626 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 417054 0 417110 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 419538 0 419594 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 225786 0 225842 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 240690 0 240746 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 268014 0 268070 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 272982 0 273038 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 277950 0 278006 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 282918 0 282974 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 292854 0 292910 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 295338 0 295394 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 300306 0 300362 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 310242 0 310298 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 317694 0 317750 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 322662 0 322718 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 325146 0 325202 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 327630 0 327686 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 337566 0 337622 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 342534 0 342590 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 345018 0 345074 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 347502 0 347558 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 349986 0 350042 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 353298 0 353354 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 355782 0 355838 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 358266 0 358322 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 360750 0 360806 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 365718 0 365774 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 368202 0 368258 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 370686 0 370742 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 373170 0 373226 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 375654 0 375710 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 378138 0 378194 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 380622 0 380678 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 383106 0 383162 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 385590 0 385646 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 388074 0 388130 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 390558 0 390614 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 393042 0 393098 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 395526 0 395582 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 398010 0 398066 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 400494 0 400550 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 402978 0 403034 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 405462 0 405518 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 407946 0 408002 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 410430 0 410486 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 412914 0 412970 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 415398 0 415454 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 417882 0 417938 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 420366 0 420422 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 144642 0 144698 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 152094 0 152150 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 196806 0 196862 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 199290 0 199346 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 204258 0 204314 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 224130 0 224186 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 226614 0 226670 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 229098 0 229154 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 234066 0 234122 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 239034 0 239090 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 246486 0 246542 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 248970 0 249026 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 256422 0 256478 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 261390 0 261446 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 263874 0 263930 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 266358 0 266414 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 273810 0 273866 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 281262 0 281318 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 283746 0 283802 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 288714 0 288770 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 291198 0 291254 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 296166 0 296222 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 298650 0 298706 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 301134 0 301190 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 303618 0 303674 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 306102 0 306158 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 308586 0 308642 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 316038 0 316094 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 318522 0 318578 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 321006 0 321062 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 323490 0 323546 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 325974 0 326030 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 330942 0 330998 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 333426 0 333482 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 335910 0 335966 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 338394 0 338450 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 340878 0 340934 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 343362 0 343418 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 348330 0 348386 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 350814 0 350870 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 356610 0 356666 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 359094 0 359150 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 361578 0 361634 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 364062 0 364118 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 366546 0 366602 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 369030 0 369086 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 371514 0 371570 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 373998 0 374054 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 378966 0 379022 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 381450 0 381506 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 383934 0 383990 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 386418 0 386474 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 388902 0 388958 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 396354 0 396410 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 398838 0 398894 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 403806 0 403862 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 406290 0 406346 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 408774 0 408830 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 411258 0 411314 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 413742 0 413798 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 416226 0 416282 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 418710 0 418766 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 277122 0 277178 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 289542 0 289598 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 292026 0 292082 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 301962 0 302018 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 304446 0 304502 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 309414 0 309470 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 319350 0 319406 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 324318 0 324374 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 326802 0 326858 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 329286 0 329342 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 331770 0 331826 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 334254 0 334310 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 336738 0 336794 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 339222 0 339278 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 341706 0 341762 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 344190 0 344246 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 346674 0 346730 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 557648 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 557648 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 16302 0 16358 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 560000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 478083166
string GDS_FILE /home/htamas/progs/trainable-nn-v3/openlane/trainable_nn/runs/22_09_13_01_49/results/signoff/trainable_nn.magic.gds
string GDS_START 1973292
<< end >>

